##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Mon Mar 10 20:20:02 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 758.0000 BY 757.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 279.7500 1.0000 280.2500 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 159.0500 0.0000 159.5500 1.0000 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 161.4500 0.0000 161.9500 1.0000 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 163.8500 0.0000 164.3500 1.0000 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 166.2500 0.0000 166.7500 1.0000 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 168.6500 0.0000 169.1500 1.0000 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 171.0500 0.0000 171.5500 1.0000 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 173.4500 0.0000 173.9500 1.0000 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 175.8500 0.0000 176.3500 1.0000 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 178.2500 0.0000 178.7500 1.0000 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 180.6500 0.0000 181.1500 1.0000 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 183.0500 0.0000 183.5500 1.0000 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 185.4500 0.0000 185.9500 1.0000 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 187.8500 0.0000 188.3500 1.0000 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 190.2500 0.0000 190.7500 1.0000 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 192.6500 0.0000 193.1500 1.0000 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 195.0500 0.0000 195.5500 1.0000 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 197.4500 0.0000 197.9500 1.0000 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 199.8500 0.0000 200.3500 1.0000 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 202.2500 0.0000 202.7500 1.0000 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 204.6500 0.0000 205.1500 1.0000 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 207.0500 0.0000 207.5500 1.0000 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 209.4500 0.0000 209.9500 1.0000 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 211.8500 0.0000 212.3500 1.0000 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 214.2500 0.0000 214.7500 1.0000 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 435.7500 1.0000 436.2500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 433.3500 1.0000 433.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 430.9500 1.0000 431.4500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 428.5500 1.0000 429.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 426.1500 1.0000 426.6500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 423.7500 1.0000 424.2500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 421.3500 1.0000 421.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 418.9500 1.0000 419.4500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 416.5500 1.0000 417.0500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 414.1500 1.0000 414.6500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 411.7500 1.0000 412.2500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 409.3500 1.0000 409.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 406.9500 1.0000 407.4500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 404.5500 1.0000 405.0500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 402.1500 1.0000 402.6500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 399.7500 1.0000 400.2500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 397.3500 1.0000 397.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 394.9500 1.0000 395.4500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 392.5500 1.0000 393.0500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 390.1500 1.0000 390.6500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 387.7500 1.0000 388.2500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 385.3500 1.0000 385.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 382.9500 1.0000 383.4500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 380.5500 1.0000 381.0500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 378.1500 1.0000 378.6500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 375.7500 1.0000 376.2500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 373.3500 1.0000 373.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 370.9500 1.0000 371.4500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 368.5500 1.0000 369.0500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 366.1500 1.0000 366.6500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 363.7500 1.0000 364.2500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 361.3500 1.0000 361.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 358.9500 1.0000 359.4500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 356.5500 1.0000 357.0500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 354.1500 1.0000 354.6500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 351.7500 1.0000 352.2500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 349.3500 1.0000 349.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 346.9500 1.0000 347.4500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 344.5500 1.0000 345.0500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 342.1500 1.0000 342.6500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 339.7500 1.0000 340.2500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 337.3500 1.0000 337.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 334.9500 1.0000 335.4500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 332.5500 1.0000 333.0500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 330.1500 1.0000 330.6500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 327.7500 1.0000 328.2500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 325.3500 1.0000 325.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 322.9500 1.0000 323.4500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 320.5500 1.0000 321.0500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 318.1500 1.0000 318.6500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 315.7500 1.0000 316.2500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 313.3500 1.0000 313.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 310.9500 1.0000 311.4500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 308.5500 1.0000 309.0500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 306.1500 1.0000 306.6500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 303.7500 1.0000 304.2500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 301.3500 1.0000 301.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 298.9500 1.0000 299.4500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 296.5500 1.0000 297.0500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 294.1500 1.0000 294.6500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 291.7500 1.0000 292.2500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 289.3500 1.0000 289.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 286.9500 1.0000 287.4500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 284.5500 1.0000 285.0500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 216.6500 0.0000 217.1500 1.0000 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 219.0500 0.0000 219.5500 1.0000 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 221.4500 0.0000 221.9500 1.0000 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 223.8500 0.0000 224.3500 1.0000 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 226.2500 0.0000 226.7500 1.0000 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 228.6500 0.0000 229.1500 1.0000 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 231.0500 0.0000 231.5500 1.0000 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 233.4500 0.0000 233.9500 1.0000 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 235.8500 0.0000 236.3500 1.0000 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 238.2500 0.0000 238.7500 1.0000 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 240.6500 0.0000 241.1500 1.0000 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 243.0500 0.0000 243.5500 1.0000 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 245.4500 0.0000 245.9500 1.0000 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 247.8500 0.0000 248.3500 1.0000 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 250.2500 0.0000 250.7500 1.0000 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 252.6500 0.0000 253.1500 1.0000 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 255.0500 0.0000 255.5500 1.0000 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 257.4500 0.0000 257.9500 1.0000 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 259.8500 0.0000 260.3500 1.0000 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 262.2500 0.0000 262.7500 1.0000 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 264.6500 0.0000 265.1500 1.0000 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 267.0500 0.0000 267.5500 1.0000 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 269.4500 0.0000 269.9500 1.0000 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 271.8500 0.0000 272.3500 1.0000 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 274.2500 0.0000 274.7500 1.0000 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 276.6500 0.0000 277.1500 1.0000 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 279.0500 0.0000 279.5500 1.0000 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 281.4500 0.0000 281.9500 1.0000 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 283.8500 0.0000 284.3500 1.0000 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 286.2500 0.0000 286.7500 1.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 288.6500 0.0000 289.1500 1.0000 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 291.0500 0.0000 291.5500 1.0000 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 293.4500 0.0000 293.9500 1.0000 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 295.8500 0.0000 296.3500 1.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 298.2500 0.0000 298.7500 1.0000 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 300.6500 0.0000 301.1500 1.0000 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 303.0500 0.0000 303.5500 1.0000 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 305.4500 0.0000 305.9500 1.0000 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 307.8500 0.0000 308.3500 1.0000 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 310.2500 0.0000 310.7500 1.0000 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 312.6500 0.0000 313.1500 1.0000 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 315.0500 0.0000 315.5500 1.0000 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 317.4500 0.0000 317.9500 1.0000 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 319.8500 0.0000 320.3500 1.0000 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 322.2500 0.0000 322.7500 1.0000 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 324.6500 0.0000 325.1500 1.0000 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 327.0500 0.0000 327.5500 1.0000 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 329.4500 0.0000 329.9500 1.0000 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 331.8500 0.0000 332.3500 1.0000 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 334.2500 0.0000 334.7500 1.0000 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 336.6500 0.0000 337.1500 1.0000 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 339.0500 0.0000 339.5500 1.0000 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 341.4500 0.0000 341.9500 1.0000 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 343.8500 0.0000 344.3500 1.0000 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 346.2500 0.0000 346.7500 1.0000 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 348.6500 0.0000 349.1500 1.0000 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 351.0500 0.0000 351.5500 1.0000 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 353.4500 0.0000 353.9500 1.0000 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 355.8500 0.0000 356.3500 1.0000 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 358.2500 0.0000 358.7500 1.0000 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 360.6500 0.0000 361.1500 1.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 363.0500 0.0000 363.5500 1.0000 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 365.4500 0.0000 365.9500 1.0000 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 367.8500 0.0000 368.3500 1.0000 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 370.2500 0.0000 370.7500 1.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 372.6500 0.0000 373.1500 1.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 375.0500 0.0000 375.5500 1.0000 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 377.4500 0.0000 377.9500 1.0000 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 379.8500 0.0000 380.3500 1.0000 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 382.2500 0.0000 382.7500 1.0000 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 384.6500 0.0000 385.1500 1.0000 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 387.0500 0.0000 387.5500 1.0000 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 389.4500 0.0000 389.9500 1.0000 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 391.8500 0.0000 392.3500 1.0000 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 394.2500 0.0000 394.7500 1.0000 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 396.6500 0.0000 397.1500 1.0000 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 399.0500 0.0000 399.5500 1.0000 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 401.4500 0.0000 401.9500 1.0000 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 403.8500 0.0000 404.3500 1.0000 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 406.2500 0.0000 406.7500 1.0000 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 408.6500 0.0000 409.1500 1.0000 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 411.0500 0.0000 411.5500 1.0000 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 413.4500 0.0000 413.9500 1.0000 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 415.8500 0.0000 416.3500 1.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 418.2500 0.0000 418.7500 1.0000 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 420.6500 0.0000 421.1500 1.0000 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 423.0500 0.0000 423.5500 1.0000 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 425.4500 0.0000 425.9500 1.0000 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 427.8500 0.0000 428.3500 1.0000 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 430.2500 0.0000 430.7500 1.0000 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 432.6500 0.0000 433.1500 1.0000 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 435.0500 0.0000 435.5500 1.0000 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 437.4500 0.0000 437.9500 1.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 439.8500 0.0000 440.3500 1.0000 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 442.2500 0.0000 442.7500 1.0000 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 444.6500 0.0000 445.1500 1.0000 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 447.0500 0.0000 447.5500 1.0000 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 449.4500 0.0000 449.9500 1.0000 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 451.8500 0.0000 452.3500 1.0000 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 454.2500 0.0000 454.7500 1.0000 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 456.6500 0.0000 457.1500 1.0000 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 459.0500 0.0000 459.5500 1.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 461.4500 0.0000 461.9500 1.0000 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 463.8500 0.0000 464.3500 1.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 466.2500 0.0000 466.7500 1.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 468.6500 0.0000 469.1500 1.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 471.0500 0.0000 471.5500 1.0000 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 473.4500 0.0000 473.9500 1.0000 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 475.8500 0.0000 476.3500 1.0000 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 478.2500 0.0000 478.7500 1.0000 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 480.6500 0.0000 481.1500 1.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 483.0500 0.0000 483.5500 1.0000 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 485.4500 0.0000 485.9500 1.0000 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 487.8500 0.0000 488.3500 1.0000 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 490.2500 0.0000 490.7500 1.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 492.6500 0.0000 493.1500 1.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 495.0500 0.0000 495.5500 1.0000 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 497.4500 0.0000 497.9500 1.0000 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 499.8500 0.0000 500.3500 1.0000 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 502.2500 0.0000 502.7500 1.0000 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 504.6500 0.0000 505.1500 1.0000 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 507.0500 0.0000 507.5500 1.0000 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 509.4500 0.0000 509.9500 1.0000 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 511.8500 0.0000 512.3500 1.0000 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 514.2500 0.0000 514.7500 1.0000 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 516.6500 0.0000 517.1500 1.0000 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 519.0500 0.0000 519.5500 1.0000 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 521.4500 0.0000 521.9500 1.0000 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.8500 0.0000 524.3500 1.0000 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 526.2500 0.0000 526.7500 1.0000 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 528.6500 0.0000 529.1500 1.0000 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 531.0500 0.0000 531.5500 1.0000 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 533.4500 0.0000 533.9500 1.0000 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 535.8500 0.0000 536.3500 1.0000 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 538.2500 0.0000 538.7500 1.0000 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 540.6500 0.0000 541.1500 1.0000 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 543.0500 0.0000 543.5500 1.0000 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 545.4500 0.0000 545.9500 1.0000 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 547.8500 0.0000 548.3500 1.0000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 550.2500 0.0000 550.7500 1.0000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 552.6500 0.0000 553.1500 1.0000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 555.0500 0.0000 555.5500 1.0000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 557.4500 0.0000 557.9500 1.0000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 559.8500 0.0000 560.3500 1.0000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 562.2500 0.0000 562.7500 1.0000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 564.6500 0.0000 565.1500 1.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 567.0500 0.0000 567.5500 1.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 569.4500 0.0000 569.9500 1.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 571.8500 0.0000 572.3500 1.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 574.2500 0.0000 574.7500 1.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 576.6500 0.0000 577.1500 1.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 579.0500 0.0000 579.5500 1.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 581.4500 0.0000 581.9500 1.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 583.8500 0.0000 584.3500 1.0000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 586.2500 0.0000 586.7500 1.0000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 588.6500 0.0000 589.1500 1.0000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 591.0500 0.0000 591.5500 1.0000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 593.4500 0.0000 593.9500 1.0000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 595.8500 0.0000 596.3500 1.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 598.2500 0.0000 598.7500 1.0000 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 476.5500 1.0000 477.0500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 474.1500 1.0000 474.6500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 471.7500 1.0000 472.2500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 469.3500 1.0000 469.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 466.9500 1.0000 467.4500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 464.5500 1.0000 465.0500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 462.1500 1.0000 462.6500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 459.7500 1.0000 460.2500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 457.3500 1.0000 457.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 454.9500 1.0000 455.4500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 452.5500 1.0000 453.0500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 450.1500 1.0000 450.6500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 447.7500 1.0000 448.2500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 445.3500 1.0000 445.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 442.9500 1.0000 443.4500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 440.5500 1.0000 441.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 438.1500 1.0000 438.6500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 282.1500 1.0000 282.6500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M3 ;
      RECT 0.0000 477.2100 758.0000 757.0000 ;
      RECT 1.1600 476.3900 758.0000 477.2100 ;
      RECT 0.0000 474.8100 758.0000 476.3900 ;
      RECT 1.1600 473.9900 758.0000 474.8100 ;
      RECT 0.0000 472.4100 758.0000 473.9900 ;
      RECT 1.1600 471.5900 758.0000 472.4100 ;
      RECT 0.0000 470.0100 758.0000 471.5900 ;
      RECT 1.1600 469.1900 758.0000 470.0100 ;
      RECT 0.0000 467.6100 758.0000 469.1900 ;
      RECT 1.1600 466.7900 758.0000 467.6100 ;
      RECT 0.0000 465.2100 758.0000 466.7900 ;
      RECT 1.1600 464.3900 758.0000 465.2100 ;
      RECT 0.0000 462.8100 758.0000 464.3900 ;
      RECT 1.1600 461.9900 758.0000 462.8100 ;
      RECT 0.0000 460.4100 758.0000 461.9900 ;
      RECT 1.1600 459.5900 758.0000 460.4100 ;
      RECT 0.0000 458.0100 758.0000 459.5900 ;
      RECT 1.1600 457.1900 758.0000 458.0100 ;
      RECT 0.0000 455.6100 758.0000 457.1900 ;
      RECT 1.1600 454.7900 758.0000 455.6100 ;
      RECT 0.0000 453.2100 758.0000 454.7900 ;
      RECT 1.1600 452.3900 758.0000 453.2100 ;
      RECT 0.0000 450.8100 758.0000 452.3900 ;
      RECT 1.1600 449.9900 758.0000 450.8100 ;
      RECT 0.0000 448.4100 758.0000 449.9900 ;
      RECT 1.1600 447.5900 758.0000 448.4100 ;
      RECT 0.0000 446.0100 758.0000 447.5900 ;
      RECT 1.1600 445.1900 758.0000 446.0100 ;
      RECT 0.0000 443.6100 758.0000 445.1900 ;
      RECT 1.1600 442.7900 758.0000 443.6100 ;
      RECT 0.0000 441.2100 758.0000 442.7900 ;
      RECT 1.1600 440.3900 758.0000 441.2100 ;
      RECT 0.0000 438.8100 758.0000 440.3900 ;
      RECT 1.1600 437.9900 758.0000 438.8100 ;
      RECT 0.0000 436.4100 758.0000 437.9900 ;
      RECT 1.1600 435.5900 758.0000 436.4100 ;
      RECT 0.0000 434.0100 758.0000 435.5900 ;
      RECT 1.1600 433.1900 758.0000 434.0100 ;
      RECT 0.0000 431.6100 758.0000 433.1900 ;
      RECT 1.1600 430.7900 758.0000 431.6100 ;
      RECT 0.0000 429.2100 758.0000 430.7900 ;
      RECT 1.1600 428.3900 758.0000 429.2100 ;
      RECT 0.0000 426.8100 758.0000 428.3900 ;
      RECT 1.1600 425.9900 758.0000 426.8100 ;
      RECT 0.0000 424.4100 758.0000 425.9900 ;
      RECT 1.1600 423.5900 758.0000 424.4100 ;
      RECT 0.0000 422.0100 758.0000 423.5900 ;
      RECT 1.1600 421.1900 758.0000 422.0100 ;
      RECT 0.0000 419.6100 758.0000 421.1900 ;
      RECT 1.1600 418.7900 758.0000 419.6100 ;
      RECT 0.0000 417.2100 758.0000 418.7900 ;
      RECT 1.1600 416.3900 758.0000 417.2100 ;
      RECT 0.0000 414.8100 758.0000 416.3900 ;
      RECT 1.1600 413.9900 758.0000 414.8100 ;
      RECT 0.0000 412.4100 758.0000 413.9900 ;
      RECT 1.1600 411.5900 758.0000 412.4100 ;
      RECT 0.0000 410.0100 758.0000 411.5900 ;
      RECT 1.1600 409.1900 758.0000 410.0100 ;
      RECT 0.0000 407.6100 758.0000 409.1900 ;
      RECT 1.1600 406.7900 758.0000 407.6100 ;
      RECT 0.0000 405.2100 758.0000 406.7900 ;
      RECT 1.1600 404.3900 758.0000 405.2100 ;
      RECT 0.0000 402.8100 758.0000 404.3900 ;
      RECT 1.1600 401.9900 758.0000 402.8100 ;
      RECT 0.0000 400.4100 758.0000 401.9900 ;
      RECT 1.1600 399.5900 758.0000 400.4100 ;
      RECT 0.0000 398.0100 758.0000 399.5900 ;
      RECT 1.1600 397.1900 758.0000 398.0100 ;
      RECT 0.0000 395.6100 758.0000 397.1900 ;
      RECT 1.1600 394.7900 758.0000 395.6100 ;
      RECT 0.0000 393.2100 758.0000 394.7900 ;
      RECT 1.1600 392.3900 758.0000 393.2100 ;
      RECT 0.0000 390.8100 758.0000 392.3900 ;
      RECT 1.1600 389.9900 758.0000 390.8100 ;
      RECT 0.0000 388.4100 758.0000 389.9900 ;
      RECT 1.1600 387.5900 758.0000 388.4100 ;
      RECT 0.0000 386.0100 758.0000 387.5900 ;
      RECT 1.1600 385.1900 758.0000 386.0100 ;
      RECT 0.0000 383.6100 758.0000 385.1900 ;
      RECT 1.1600 382.7900 758.0000 383.6100 ;
      RECT 0.0000 381.2100 758.0000 382.7900 ;
      RECT 1.1600 380.3900 758.0000 381.2100 ;
      RECT 0.0000 378.8100 758.0000 380.3900 ;
      RECT 1.1600 377.9900 758.0000 378.8100 ;
      RECT 0.0000 376.4100 758.0000 377.9900 ;
      RECT 1.1600 375.5900 758.0000 376.4100 ;
      RECT 0.0000 374.0100 758.0000 375.5900 ;
      RECT 1.1600 373.1900 758.0000 374.0100 ;
      RECT 0.0000 371.6100 758.0000 373.1900 ;
      RECT 1.1600 370.7900 758.0000 371.6100 ;
      RECT 0.0000 369.2100 758.0000 370.7900 ;
      RECT 1.1600 368.3900 758.0000 369.2100 ;
      RECT 0.0000 366.8100 758.0000 368.3900 ;
      RECT 1.1600 365.9900 758.0000 366.8100 ;
      RECT 0.0000 364.4100 758.0000 365.9900 ;
      RECT 1.1600 363.5900 758.0000 364.4100 ;
      RECT 0.0000 362.0100 758.0000 363.5900 ;
      RECT 1.1600 361.1900 758.0000 362.0100 ;
      RECT 0.0000 359.6100 758.0000 361.1900 ;
      RECT 1.1600 358.7900 758.0000 359.6100 ;
      RECT 0.0000 357.2100 758.0000 358.7900 ;
      RECT 1.1600 356.3900 758.0000 357.2100 ;
      RECT 0.0000 354.8100 758.0000 356.3900 ;
      RECT 1.1600 353.9900 758.0000 354.8100 ;
      RECT 0.0000 352.4100 758.0000 353.9900 ;
      RECT 1.1600 351.5900 758.0000 352.4100 ;
      RECT 0.0000 350.0100 758.0000 351.5900 ;
      RECT 1.1600 349.1900 758.0000 350.0100 ;
      RECT 0.0000 347.6100 758.0000 349.1900 ;
      RECT 1.1600 346.7900 758.0000 347.6100 ;
      RECT 0.0000 345.2100 758.0000 346.7900 ;
      RECT 1.1600 344.3900 758.0000 345.2100 ;
      RECT 0.0000 342.8100 758.0000 344.3900 ;
      RECT 1.1600 341.9900 758.0000 342.8100 ;
      RECT 0.0000 340.4100 758.0000 341.9900 ;
      RECT 1.1600 339.5900 758.0000 340.4100 ;
      RECT 0.0000 338.0100 758.0000 339.5900 ;
      RECT 1.1600 337.1900 758.0000 338.0100 ;
      RECT 0.0000 335.6100 758.0000 337.1900 ;
      RECT 1.1600 334.7900 758.0000 335.6100 ;
      RECT 0.0000 333.2100 758.0000 334.7900 ;
      RECT 1.1600 332.3900 758.0000 333.2100 ;
      RECT 0.0000 330.8100 758.0000 332.3900 ;
      RECT 1.1600 329.9900 758.0000 330.8100 ;
      RECT 0.0000 328.4100 758.0000 329.9900 ;
      RECT 1.1600 327.5900 758.0000 328.4100 ;
      RECT 0.0000 326.0100 758.0000 327.5900 ;
      RECT 1.1600 325.1900 758.0000 326.0100 ;
      RECT 0.0000 323.6100 758.0000 325.1900 ;
      RECT 1.1600 322.7900 758.0000 323.6100 ;
      RECT 0.0000 321.2100 758.0000 322.7900 ;
      RECT 1.1600 320.3900 758.0000 321.2100 ;
      RECT 0.0000 318.8100 758.0000 320.3900 ;
      RECT 1.1600 317.9900 758.0000 318.8100 ;
      RECT 0.0000 316.4100 758.0000 317.9900 ;
      RECT 1.1600 315.5900 758.0000 316.4100 ;
      RECT 0.0000 314.0100 758.0000 315.5900 ;
      RECT 1.1600 313.1900 758.0000 314.0100 ;
      RECT 0.0000 311.6100 758.0000 313.1900 ;
      RECT 1.1600 310.7900 758.0000 311.6100 ;
      RECT 0.0000 309.2100 758.0000 310.7900 ;
      RECT 1.1600 308.3900 758.0000 309.2100 ;
      RECT 0.0000 306.8100 758.0000 308.3900 ;
      RECT 1.1600 305.9900 758.0000 306.8100 ;
      RECT 0.0000 304.4100 758.0000 305.9900 ;
      RECT 1.1600 303.5900 758.0000 304.4100 ;
      RECT 0.0000 302.0100 758.0000 303.5900 ;
      RECT 1.1600 301.1900 758.0000 302.0100 ;
      RECT 0.0000 299.6100 758.0000 301.1900 ;
      RECT 1.1600 298.7900 758.0000 299.6100 ;
      RECT 0.0000 297.2100 758.0000 298.7900 ;
      RECT 1.1600 296.3900 758.0000 297.2100 ;
      RECT 0.0000 294.8100 758.0000 296.3900 ;
      RECT 1.1600 293.9900 758.0000 294.8100 ;
      RECT 0.0000 292.4100 758.0000 293.9900 ;
      RECT 1.1600 291.5900 758.0000 292.4100 ;
      RECT 0.0000 290.0100 758.0000 291.5900 ;
      RECT 1.1600 289.1900 758.0000 290.0100 ;
      RECT 0.0000 287.6100 758.0000 289.1900 ;
      RECT 1.1600 286.7900 758.0000 287.6100 ;
      RECT 0.0000 285.2100 758.0000 286.7900 ;
      RECT 1.1600 284.3900 758.0000 285.2100 ;
      RECT 0.0000 282.8100 758.0000 284.3900 ;
      RECT 1.1600 281.9900 758.0000 282.8100 ;
      RECT 0.0000 280.4100 758.0000 281.9900 ;
      RECT 1.1600 279.5900 758.0000 280.4100 ;
      RECT 0.0000 1.1600 758.0000 279.5900 ;
      RECT 598.9100 0.0000 758.0000 1.1600 ;
      RECT 596.5100 0.0000 598.0900 1.1600 ;
      RECT 594.1100 0.0000 595.6900 1.1600 ;
      RECT 591.7100 0.0000 593.2900 1.1600 ;
      RECT 589.3100 0.0000 590.8900 1.1600 ;
      RECT 586.9100 0.0000 588.4900 1.1600 ;
      RECT 584.5100 0.0000 586.0900 1.1600 ;
      RECT 582.1100 0.0000 583.6900 1.1600 ;
      RECT 579.7100 0.0000 581.2900 1.1600 ;
      RECT 577.3100 0.0000 578.8900 1.1600 ;
      RECT 574.9100 0.0000 576.4900 1.1600 ;
      RECT 572.5100 0.0000 574.0900 1.1600 ;
      RECT 570.1100 0.0000 571.6900 1.1600 ;
      RECT 567.7100 0.0000 569.2900 1.1600 ;
      RECT 565.3100 0.0000 566.8900 1.1600 ;
      RECT 562.9100 0.0000 564.4900 1.1600 ;
      RECT 560.5100 0.0000 562.0900 1.1600 ;
      RECT 558.1100 0.0000 559.6900 1.1600 ;
      RECT 555.7100 0.0000 557.2900 1.1600 ;
      RECT 553.3100 0.0000 554.8900 1.1600 ;
      RECT 550.9100 0.0000 552.4900 1.1600 ;
      RECT 548.5100 0.0000 550.0900 1.1600 ;
      RECT 546.1100 0.0000 547.6900 1.1600 ;
      RECT 543.7100 0.0000 545.2900 1.1600 ;
      RECT 541.3100 0.0000 542.8900 1.1600 ;
      RECT 538.9100 0.0000 540.4900 1.1600 ;
      RECT 536.5100 0.0000 538.0900 1.1600 ;
      RECT 534.1100 0.0000 535.6900 1.1600 ;
      RECT 531.7100 0.0000 533.2900 1.1600 ;
      RECT 529.3100 0.0000 530.8900 1.1600 ;
      RECT 526.9100 0.0000 528.4900 1.1600 ;
      RECT 524.5100 0.0000 526.0900 1.1600 ;
      RECT 522.1100 0.0000 523.6900 1.1600 ;
      RECT 519.7100 0.0000 521.2900 1.1600 ;
      RECT 517.3100 0.0000 518.8900 1.1600 ;
      RECT 514.9100 0.0000 516.4900 1.1600 ;
      RECT 512.5100 0.0000 514.0900 1.1600 ;
      RECT 510.1100 0.0000 511.6900 1.1600 ;
      RECT 507.7100 0.0000 509.2900 1.1600 ;
      RECT 505.3100 0.0000 506.8900 1.1600 ;
      RECT 502.9100 0.0000 504.4900 1.1600 ;
      RECT 500.5100 0.0000 502.0900 1.1600 ;
      RECT 498.1100 0.0000 499.6900 1.1600 ;
      RECT 495.7100 0.0000 497.2900 1.1600 ;
      RECT 493.3100 0.0000 494.8900 1.1600 ;
      RECT 490.9100 0.0000 492.4900 1.1600 ;
      RECT 488.5100 0.0000 490.0900 1.1600 ;
      RECT 486.1100 0.0000 487.6900 1.1600 ;
      RECT 483.7100 0.0000 485.2900 1.1600 ;
      RECT 481.3100 0.0000 482.8900 1.1600 ;
      RECT 478.9100 0.0000 480.4900 1.1600 ;
      RECT 476.5100 0.0000 478.0900 1.1600 ;
      RECT 474.1100 0.0000 475.6900 1.1600 ;
      RECT 471.7100 0.0000 473.2900 1.1600 ;
      RECT 469.3100 0.0000 470.8900 1.1600 ;
      RECT 466.9100 0.0000 468.4900 1.1600 ;
      RECT 464.5100 0.0000 466.0900 1.1600 ;
      RECT 462.1100 0.0000 463.6900 1.1600 ;
      RECT 459.7100 0.0000 461.2900 1.1600 ;
      RECT 457.3100 0.0000 458.8900 1.1600 ;
      RECT 454.9100 0.0000 456.4900 1.1600 ;
      RECT 452.5100 0.0000 454.0900 1.1600 ;
      RECT 450.1100 0.0000 451.6900 1.1600 ;
      RECT 447.7100 0.0000 449.2900 1.1600 ;
      RECT 445.3100 0.0000 446.8900 1.1600 ;
      RECT 442.9100 0.0000 444.4900 1.1600 ;
      RECT 440.5100 0.0000 442.0900 1.1600 ;
      RECT 438.1100 0.0000 439.6900 1.1600 ;
      RECT 435.7100 0.0000 437.2900 1.1600 ;
      RECT 433.3100 0.0000 434.8900 1.1600 ;
      RECT 430.9100 0.0000 432.4900 1.1600 ;
      RECT 428.5100 0.0000 430.0900 1.1600 ;
      RECT 426.1100 0.0000 427.6900 1.1600 ;
      RECT 423.7100 0.0000 425.2900 1.1600 ;
      RECT 421.3100 0.0000 422.8900 1.1600 ;
      RECT 418.9100 0.0000 420.4900 1.1600 ;
      RECT 416.5100 0.0000 418.0900 1.1600 ;
      RECT 414.1100 0.0000 415.6900 1.1600 ;
      RECT 411.7100 0.0000 413.2900 1.1600 ;
      RECT 409.3100 0.0000 410.8900 1.1600 ;
      RECT 406.9100 0.0000 408.4900 1.1600 ;
      RECT 404.5100 0.0000 406.0900 1.1600 ;
      RECT 402.1100 0.0000 403.6900 1.1600 ;
      RECT 399.7100 0.0000 401.2900 1.1600 ;
      RECT 397.3100 0.0000 398.8900 1.1600 ;
      RECT 394.9100 0.0000 396.4900 1.1600 ;
      RECT 392.5100 0.0000 394.0900 1.1600 ;
      RECT 390.1100 0.0000 391.6900 1.1600 ;
      RECT 387.7100 0.0000 389.2900 1.1600 ;
      RECT 385.3100 0.0000 386.8900 1.1600 ;
      RECT 382.9100 0.0000 384.4900 1.1600 ;
      RECT 380.5100 0.0000 382.0900 1.1600 ;
      RECT 378.1100 0.0000 379.6900 1.1600 ;
      RECT 375.7100 0.0000 377.2900 1.1600 ;
      RECT 373.3100 0.0000 374.8900 1.1600 ;
      RECT 370.9100 0.0000 372.4900 1.1600 ;
      RECT 368.5100 0.0000 370.0900 1.1600 ;
      RECT 366.1100 0.0000 367.6900 1.1600 ;
      RECT 363.7100 0.0000 365.2900 1.1600 ;
      RECT 361.3100 0.0000 362.8900 1.1600 ;
      RECT 358.9100 0.0000 360.4900 1.1600 ;
      RECT 356.5100 0.0000 358.0900 1.1600 ;
      RECT 354.1100 0.0000 355.6900 1.1600 ;
      RECT 351.7100 0.0000 353.2900 1.1600 ;
      RECT 349.3100 0.0000 350.8900 1.1600 ;
      RECT 346.9100 0.0000 348.4900 1.1600 ;
      RECT 344.5100 0.0000 346.0900 1.1600 ;
      RECT 342.1100 0.0000 343.6900 1.1600 ;
      RECT 339.7100 0.0000 341.2900 1.1600 ;
      RECT 337.3100 0.0000 338.8900 1.1600 ;
      RECT 334.9100 0.0000 336.4900 1.1600 ;
      RECT 332.5100 0.0000 334.0900 1.1600 ;
      RECT 330.1100 0.0000 331.6900 1.1600 ;
      RECT 327.7100 0.0000 329.2900 1.1600 ;
      RECT 325.3100 0.0000 326.8900 1.1600 ;
      RECT 322.9100 0.0000 324.4900 1.1600 ;
      RECT 320.5100 0.0000 322.0900 1.1600 ;
      RECT 318.1100 0.0000 319.6900 1.1600 ;
      RECT 315.7100 0.0000 317.2900 1.1600 ;
      RECT 313.3100 0.0000 314.8900 1.1600 ;
      RECT 310.9100 0.0000 312.4900 1.1600 ;
      RECT 308.5100 0.0000 310.0900 1.1600 ;
      RECT 306.1100 0.0000 307.6900 1.1600 ;
      RECT 303.7100 0.0000 305.2900 1.1600 ;
      RECT 301.3100 0.0000 302.8900 1.1600 ;
      RECT 298.9100 0.0000 300.4900 1.1600 ;
      RECT 296.5100 0.0000 298.0900 1.1600 ;
      RECT 294.1100 0.0000 295.6900 1.1600 ;
      RECT 291.7100 0.0000 293.2900 1.1600 ;
      RECT 289.3100 0.0000 290.8900 1.1600 ;
      RECT 286.9100 0.0000 288.4900 1.1600 ;
      RECT 284.5100 0.0000 286.0900 1.1600 ;
      RECT 282.1100 0.0000 283.6900 1.1600 ;
      RECT 279.7100 0.0000 281.2900 1.1600 ;
      RECT 277.3100 0.0000 278.8900 1.1600 ;
      RECT 274.9100 0.0000 276.4900 1.1600 ;
      RECT 272.5100 0.0000 274.0900 1.1600 ;
      RECT 270.1100 0.0000 271.6900 1.1600 ;
      RECT 267.7100 0.0000 269.2900 1.1600 ;
      RECT 265.3100 0.0000 266.8900 1.1600 ;
      RECT 262.9100 0.0000 264.4900 1.1600 ;
      RECT 260.5100 0.0000 262.0900 1.1600 ;
      RECT 258.1100 0.0000 259.6900 1.1600 ;
      RECT 255.7100 0.0000 257.2900 1.1600 ;
      RECT 253.3100 0.0000 254.8900 1.1600 ;
      RECT 250.9100 0.0000 252.4900 1.1600 ;
      RECT 248.5100 0.0000 250.0900 1.1600 ;
      RECT 246.1100 0.0000 247.6900 1.1600 ;
      RECT 243.7100 0.0000 245.2900 1.1600 ;
      RECT 241.3100 0.0000 242.8900 1.1600 ;
      RECT 238.9100 0.0000 240.4900 1.1600 ;
      RECT 236.5100 0.0000 238.0900 1.1600 ;
      RECT 234.1100 0.0000 235.6900 1.1600 ;
      RECT 231.7100 0.0000 233.2900 1.1600 ;
      RECT 229.3100 0.0000 230.8900 1.1600 ;
      RECT 226.9100 0.0000 228.4900 1.1600 ;
      RECT 224.5100 0.0000 226.0900 1.1600 ;
      RECT 222.1100 0.0000 223.6900 1.1600 ;
      RECT 219.7100 0.0000 221.2900 1.1600 ;
      RECT 217.3100 0.0000 218.8900 1.1600 ;
      RECT 214.9100 0.0000 216.4900 1.1600 ;
      RECT 212.5100 0.0000 214.0900 1.1600 ;
      RECT 210.1100 0.0000 211.6900 1.1600 ;
      RECT 207.7100 0.0000 209.2900 1.1600 ;
      RECT 205.3100 0.0000 206.8900 1.1600 ;
      RECT 202.9100 0.0000 204.4900 1.1600 ;
      RECT 200.5100 0.0000 202.0900 1.1600 ;
      RECT 198.1100 0.0000 199.6900 1.1600 ;
      RECT 195.7100 0.0000 197.2900 1.1600 ;
      RECT 193.3100 0.0000 194.8900 1.1600 ;
      RECT 190.9100 0.0000 192.4900 1.1600 ;
      RECT 188.5100 0.0000 190.0900 1.1600 ;
      RECT 186.1100 0.0000 187.6900 1.1600 ;
      RECT 183.7100 0.0000 185.2900 1.1600 ;
      RECT 181.3100 0.0000 182.8900 1.1600 ;
      RECT 178.9100 0.0000 180.4900 1.1600 ;
      RECT 176.5100 0.0000 178.0900 1.1600 ;
      RECT 174.1100 0.0000 175.6900 1.1600 ;
      RECT 171.7100 0.0000 173.2900 1.1600 ;
      RECT 169.3100 0.0000 170.8900 1.1600 ;
      RECT 166.9100 0.0000 168.4900 1.1600 ;
      RECT 164.5100 0.0000 166.0900 1.1600 ;
      RECT 162.1100 0.0000 163.6900 1.1600 ;
      RECT 159.7100 0.0000 161.2900 1.1600 ;
      RECT 0.0000 0.0000 158.8900 1.1600 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 758.0000 757.0000 ;
  END
END core

END LIBRARY
