##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sun Feb 16 19:53:55 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO add
  CLASS BLOCK ;
  SIZE 40.8000 BY 38.0000 ;
  FOREIGN add 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.4500 37.4800 18.5500 38.0000 ;
    END
  END clk
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 40.2800 14.9500 40.8000 15.0500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0500 0.0000 29.1500 0.5200 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 40.2800 19.3500 40.8000 19.4500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 40.2800 25.7500 40.8000 25.8500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.0500 37.4800 29.1500 38.0000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 40.2800 18.5500 40.8000 18.6500 ;
    END
  END out[0]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.0500 0.0000 16.1500 0.5200 ;
    END
  END x[3]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.3500 0.5200 23.4500 ;
    END
  END x[2]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.0500 37.4800 14.1500 38.0000 ;
    END
  END x[1]
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.1500 0.5200 18.2500 ;
    END
  END x[0]
  PIN y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 16.0500 0.0000 16.1500 0.5200 ;
    END
  END y[3]
  PIN y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.7500 0.5200 19.8500 ;
    END
  END y[2]
  PIN y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 14.2500 37.4800 14.3500 38.0000 ;
    END
  END y[1]
  PIN y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.1500 0.5200 16.2500 ;
    END
  END y[0]
  PIN z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.0500 0.0000 14.1500 0.5200 ;
    END
  END z[3]
  PIN z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.6500 37.4800 19.7500 38.0000 ;
    END
  END z[2]
  PIN z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 37.4800 18.1500 38.0000 ;
    END
  END z[1]
  PIN z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.0500 0.0000 18.1500 0.5200 ;
    END
  END z[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 40.8000 38.0000 ;
    LAYER M2 ;
      RECT 29.2500 37.3800 40.8000 38.0000 ;
      RECT 19.8500 37.3800 28.9500 38.0000 ;
      RECT 18.6500 37.3800 19.5500 38.0000 ;
      RECT 18.2500 37.3800 18.3500 38.0000 ;
      RECT 14.2500 37.3800 17.9500 38.0000 ;
      RECT 0.0000 37.3800 13.9500 38.0000 ;
      RECT 0.0000 0.6200 40.8000 37.3800 ;
      RECT 29.2500 0.0000 40.8000 0.6200 ;
      RECT 18.2500 0.0000 28.9500 0.6200 ;
      RECT 16.2500 0.0000 17.9500 0.6200 ;
      RECT 14.2500 0.0000 15.9500 0.6200 ;
      RECT 0.0000 0.0000 13.9500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 25.9500 40.8000 38.0000 ;
      RECT 0.0000 25.6500 40.1800 25.9500 ;
      RECT 0.0000 23.5500 40.8000 25.6500 ;
      RECT 0.6200 23.2500 40.8000 23.5500 ;
      RECT 0.0000 19.9500 40.8000 23.2500 ;
      RECT 0.6200 19.6500 40.8000 19.9500 ;
      RECT 0.0000 19.5500 40.8000 19.6500 ;
      RECT 0.0000 19.2500 40.1800 19.5500 ;
      RECT 0.0000 18.7500 40.8000 19.2500 ;
      RECT 0.0000 18.4500 40.1800 18.7500 ;
      RECT 0.0000 18.3500 40.8000 18.4500 ;
      RECT 0.6200 18.0500 40.8000 18.3500 ;
      RECT 0.0000 16.3500 40.8000 18.0500 ;
      RECT 0.6200 16.0500 40.8000 16.3500 ;
      RECT 0.0000 15.1500 40.8000 16.0500 ;
      RECT 0.0000 14.8500 40.1800 15.1500 ;
      RECT 0.0000 0.0000 40.8000 14.8500 ;
    LAYER M4 ;
      RECT 14.4500 37.3800 40.8000 38.0000 ;
      RECT 0.0000 37.3800 14.1500 38.0000 ;
      RECT 0.0000 0.6200 40.8000 37.3800 ;
      RECT 16.2500 0.0000 40.8000 0.6200 ;
      RECT 0.0000 0.0000 15.9500 0.6200 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 40.8000 38.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 40.8000 38.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 40.8000 38.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 40.8000 38.0000 ;
  END
END add

END LIBRARY
