##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar 21 21:15:34 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 346.4000 BY 344.8000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.9500 0.6000 20.0500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.4500 0.0000 122.5500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.2500 0.0000 123.3500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0500 0.0000 124.1500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 0.0000 124.9500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.6500 0.0000 125.7500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.4500 0.0000 126.5500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.2500 0.0000 127.3500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.0500 0.0000 128.1500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 0.0000 128.9500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.6500 0.0000 129.7500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.4500 0.0000 130.5500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.2500 0.0000 131.3500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.0500 0.0000 132.1500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 0.0000 132.9500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.6500 0.0000 133.7500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.4500 0.0000 134.5500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.2500 0.0000 135.3500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.0500 0.0000 136.1500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 0.0000 136.9500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.6500 0.0000 137.7500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.4500 0.0000 138.5500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.2500 0.0000 139.3500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.0500 0.0000 140.1500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 0.0000 140.9500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.6500 0.0000 141.7500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.4500 0.0000 142.5500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.2500 0.0000 143.3500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.0500 0.0000 144.1500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 0.0000 144.9500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.6500 0.0000 145.7500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.4500 0.0000 146.5500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.2500 0.0000 147.3500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.0500 0.0000 148.1500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 0.0000 148.9500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.6500 0.0000 149.7500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.4500 0.0000 150.5500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.2500 0.0000 151.3500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.0500 0.0000 152.1500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 0.0000 152.9500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.6500 0.0000 153.7500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.4500 0.0000 154.5500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.2500 0.0000 155.3500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.0500 0.0000 156.1500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 0.0000 156.9500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.6500 0.0000 157.7500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.4500 0.0000 158.5500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.2500 0.0000 159.3500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.0500 0.0000 160.1500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 0.0000 160.9500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.6500 0.0000 161.7500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.4500 0.0000 162.5500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.2500 0.0000 163.3500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.0500 0.0000 164.1500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 0.0000 164.9500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.6500 0.0000 165.7500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.4500 0.0000 166.5500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.2500 0.0000 167.3500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.0500 0.0000 168.1500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 0.0000 168.9500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.6500 0.0000 169.7500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.4500 0.0000 170.5500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.2500 0.0000 171.3500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.0500 0.0000 172.1500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.8500 0.0000 172.9500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.6500 0.0000 173.7500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.4500 0.0000 174.5500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.2500 0.0000 175.3500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.0500 0.0000 176.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.8500 0.0000 176.9500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.6500 0.0000 177.7500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.4500 0.0000 178.5500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.2500 0.0000 179.3500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.0500 0.0000 180.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.8500 0.0000 180.9500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.6500 0.0000 181.7500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.4500 0.0000 182.5500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.2500 0.0000 183.3500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.0500 0.0000 184.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.8500 0.0000 184.9500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.6500 0.0000 185.7500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.4500 0.0000 186.5500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.2500 0.0000 187.3500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.0500 0.0000 188.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.8500 0.0000 188.9500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.6500 0.0000 189.7500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.4500 0.0000 190.5500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.2500 0.0000 191.3500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.0500 0.0000 192.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.8500 0.0000 192.9500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.6500 0.0000 193.7500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.4500 0.0000 194.5500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.2500 0.0000 195.3500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.0500 0.0000 196.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.8500 0.0000 196.9500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.6500 0.0000 197.7500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.4500 0.0000 198.5500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.2500 0.0000 199.3500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.0500 0.0000 200.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.8500 0.0000 200.9500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.6500 0.0000 201.7500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.4500 0.0000 202.5500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.2500 0.0000 203.3500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.0500 0.0000 204.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.8500 0.0000 204.9500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.6500 0.0000 205.7500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.4500 0.0000 206.5500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.2500 0.0000 207.3500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.0500 0.0000 208.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.8500 0.0000 208.9500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.6500 0.0000 209.7500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.4500 0.0000 210.5500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.2500 0.0000 211.3500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.0500 0.0000 212.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.8500 0.0000 212.9500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.6500 0.0000 213.7500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.4500 0.0000 214.5500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.2500 0.0000 215.3500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.0500 0.0000 216.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.8500 0.0000 216.9500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.6500 0.0000 217.7500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.4500 0.0000 218.5500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.2500 0.0000 219.3500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.0500 0.0000 220.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.8500 0.0000 220.9500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.6500 0.0000 221.7500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.4500 0.0000 222.5500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.2500 0.0000 223.3500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.0500 0.0000 224.1500 0.6000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.4500 344.2000 122.5500 344.8000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.2500 344.2000 123.3500 344.8000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0500 344.2000 124.1500 344.8000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.8500 344.2000 124.9500 344.8000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.6500 344.2000 125.7500 344.8000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.4500 344.2000 126.5500 344.8000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.2500 344.2000 127.3500 344.8000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.0500 344.2000 128.1500 344.8000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.8500 344.2000 128.9500 344.8000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.6500 344.2000 129.7500 344.8000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.4500 344.2000 130.5500 344.8000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.2500 344.2000 131.3500 344.8000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.0500 344.2000 132.1500 344.8000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.8500 344.2000 132.9500 344.8000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.6500 344.2000 133.7500 344.8000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.4500 344.2000 134.5500 344.8000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.2500 344.2000 135.3500 344.8000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.0500 344.2000 136.1500 344.8000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.8500 344.2000 136.9500 344.8000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.6500 344.2000 137.7500 344.8000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.4500 344.2000 138.5500 344.8000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.2500 344.2000 139.3500 344.8000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.0500 344.2000 140.1500 344.8000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.8500 344.2000 140.9500 344.8000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.6500 344.2000 141.7500 344.8000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.4500 344.2000 142.5500 344.8000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.2500 344.2000 143.3500 344.8000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.0500 344.2000 144.1500 344.8000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.8500 344.2000 144.9500 344.8000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.6500 344.2000 145.7500 344.8000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.4500 344.2000 146.5500 344.8000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.2500 344.2000 147.3500 344.8000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.0500 344.2000 148.1500 344.8000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.8500 344.2000 148.9500 344.8000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.6500 344.2000 149.7500 344.8000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.4500 344.2000 150.5500 344.8000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.2500 344.2000 151.3500 344.8000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.0500 344.2000 152.1500 344.8000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.8500 344.2000 152.9500 344.8000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.6500 344.2000 153.7500 344.8000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.4500 344.2000 154.5500 344.8000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.2500 344.2000 155.3500 344.8000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.0500 344.2000 156.1500 344.8000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.8500 344.2000 156.9500 344.8000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.6500 344.2000 157.7500 344.8000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.4500 344.2000 158.5500 344.8000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.2500 344.2000 159.3500 344.8000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.0500 344.2000 160.1500 344.8000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.8500 344.2000 160.9500 344.8000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.6500 344.2000 161.7500 344.8000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.4500 344.2000 162.5500 344.8000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.2500 344.2000 163.3500 344.8000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.0500 344.2000 164.1500 344.8000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 344.2000 164.9500 344.8000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.6500 344.2000 165.7500 344.8000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.4500 344.2000 166.5500 344.8000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.2500 344.2000 167.3500 344.8000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.0500 344.2000 168.1500 344.8000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.8500 344.2000 168.9500 344.8000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.6500 344.2000 169.7500 344.8000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.4500 344.2000 170.5500 344.8000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.2500 344.2000 171.3500 344.8000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.0500 344.2000 172.1500 344.8000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.8500 344.2000 172.9500 344.8000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.6500 344.2000 173.7500 344.8000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.4500 344.2000 174.5500 344.8000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.2500 344.2000 175.3500 344.8000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.0500 344.2000 176.1500 344.8000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.8500 344.2000 176.9500 344.8000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.6500 344.2000 177.7500 344.8000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.4500 344.2000 178.5500 344.8000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.2500 344.2000 179.3500 344.8000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.0500 344.2000 180.1500 344.8000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.8500 344.2000 180.9500 344.8000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.6500 344.2000 181.7500 344.8000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.4500 344.2000 182.5500 344.8000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.2500 344.2000 183.3500 344.8000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.0500 344.2000 184.1500 344.8000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.8500 344.2000 184.9500 344.8000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.6500 344.2000 185.7500 344.8000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.4500 344.2000 186.5500 344.8000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.2500 344.2000 187.3500 344.8000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.0500 344.2000 188.1500 344.8000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.8500 344.2000 188.9500 344.8000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.6500 344.2000 189.7500 344.8000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.4500 344.2000 190.5500 344.8000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.2500 344.2000 191.3500 344.8000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.0500 344.2000 192.1500 344.8000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.8500 344.2000 192.9500 344.8000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.6500 344.2000 193.7500 344.8000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.4500 344.2000 194.5500 344.8000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.2500 344.2000 195.3500 344.8000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.0500 344.2000 196.1500 344.8000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.8500 344.2000 196.9500 344.8000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.6500 344.2000 197.7500 344.8000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.4500 344.2000 198.5500 344.8000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.2500 344.2000 199.3500 344.8000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.0500 344.2000 200.1500 344.8000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.8500 344.2000 200.9500 344.8000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.6500 344.2000 201.7500 344.8000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.4500 344.2000 202.5500 344.8000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.2500 344.2000 203.3500 344.8000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.0500 344.2000 204.1500 344.8000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.8500 344.2000 204.9500 344.8000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.6500 344.2000 205.7500 344.8000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 206.4500 344.2000 206.5500 344.8000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.2500 344.2000 207.3500 344.8000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.0500 344.2000 208.1500 344.8000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.8500 344.2000 208.9500 344.8000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.6500 344.2000 209.7500 344.8000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.4500 344.2000 210.5500 344.8000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.2500 344.2000 211.3500 344.8000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.0500 344.2000 212.1500 344.8000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.8500 344.2000 212.9500 344.8000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.6500 344.2000 213.7500 344.8000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.4500 344.2000 214.5500 344.8000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.2500 344.2000 215.3500 344.8000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.0500 344.2000 216.1500 344.8000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.8500 344.2000 216.9500 344.8000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.6500 344.2000 217.7500 344.8000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.4500 344.2000 218.5500 344.8000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.2500 344.2000 219.3500 344.8000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.0500 344.2000 220.1500 344.8000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.8500 344.2000 220.9500 344.8000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.6500 344.2000 221.7500 344.8000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.4500 344.2000 222.5500 344.8000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.2500 344.2000 223.3500 344.8000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.0500 344.2000 224.1500 344.8000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.1500 0.6000 19.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.7500 0.6000 20.8500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.3500 0.6000 18.4500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.5500 0.6000 17.6500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7500 0.6000 16.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.9500 0.6000 16.0500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 58.0000 50.0000 60.0000 294.8000 ;
        RECT 84.2650 50.0000 86.2650 294.8000 ;
        RECT 110.5300 50.0000 112.5300 294.8000 ;
        RECT 136.7950 50.0000 138.7950 294.8000 ;
        RECT 163.0600 50.0000 165.0600 294.8000 ;
        RECT 189.3250 50.0000 191.3250 294.8000 ;
        RECT 215.5900 50.0000 217.5900 294.8000 ;
        RECT 241.8550 50.0000 243.8550 294.8000 ;
        RECT 268.1200 50.0000 270.1200 294.8000 ;
        RECT 294.3850 50.0000 296.3850 294.8000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 50.0000 50.0000 52.0000 294.8000 ;
        RECT 76.2650 50.0000 78.2650 294.8000 ;
        RECT 102.5300 50.0000 104.5300 294.8000 ;
        RECT 128.7950 50.0000 130.7950 294.8000 ;
        RECT 155.0600 50.0000 157.0600 294.8000 ;
        RECT 181.3250 50.0000 183.3250 294.8000 ;
        RECT 207.5900 50.0000 209.5900 294.8000 ;
        RECT 233.8550 50.0000 235.8550 294.8000 ;
        RECT 260.1200 50.0000 262.1200 294.8000 ;
        RECT 286.3850 50.0000 288.3850 294.8000 ;
        RECT 50.0000 49.8350 52.0000 50.1650 ;
        RECT 76.2650 49.8350 78.2650 50.1650 ;
        RECT 128.7950 49.8350 130.7950 50.1650 ;
        RECT 102.5300 49.8350 104.5300 50.1650 ;
        RECT 155.0600 49.8350 157.0600 50.1650 ;
        RECT 181.3250 49.8350 183.3250 50.1650 ;
        RECT 207.5900 49.8350 209.5900 50.1650 ;
        RECT 233.8550 49.8350 235.8550 50.1650 ;
        RECT 260.1200 49.8350 262.1200 50.1650 ;
        RECT 286.3850 49.8350 288.3850 50.1650 ;
        RECT 50.0000 294.6350 52.0000 294.9650 ;
        RECT 76.2650 294.6350 78.2650 294.9650 ;
        RECT 128.7950 294.6350 130.7950 294.9650 ;
        RECT 102.5300 294.6350 104.5300 294.9650 ;
        RECT 155.0600 294.6350 157.0600 294.9650 ;
        RECT 181.3250 294.6350 183.3250 294.9650 ;
        RECT 207.5900 294.6350 209.5900 294.9650 ;
        RECT 233.8550 294.6350 235.8550 294.9650 ;
        RECT 260.1200 294.6350 262.1200 294.9650 ;
        RECT 286.3850 294.6350 288.3850 294.9650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 346.4000 344.8000 ;
    LAYER M2 ;
      RECT 224.2500 344.1000 346.4000 344.8000 ;
      RECT 223.4500 344.1000 223.9500 344.8000 ;
      RECT 222.6500 344.1000 223.1500 344.8000 ;
      RECT 221.8500 344.1000 222.3500 344.8000 ;
      RECT 221.0500 344.1000 221.5500 344.8000 ;
      RECT 220.2500 344.1000 220.7500 344.8000 ;
      RECT 219.4500 344.1000 219.9500 344.8000 ;
      RECT 218.6500 344.1000 219.1500 344.8000 ;
      RECT 217.8500 344.1000 218.3500 344.8000 ;
      RECT 217.0500 344.1000 217.5500 344.8000 ;
      RECT 216.2500 344.1000 216.7500 344.8000 ;
      RECT 215.4500 344.1000 215.9500 344.8000 ;
      RECT 214.6500 344.1000 215.1500 344.8000 ;
      RECT 213.8500 344.1000 214.3500 344.8000 ;
      RECT 213.0500 344.1000 213.5500 344.8000 ;
      RECT 212.2500 344.1000 212.7500 344.8000 ;
      RECT 211.4500 344.1000 211.9500 344.8000 ;
      RECT 210.6500 344.1000 211.1500 344.8000 ;
      RECT 209.8500 344.1000 210.3500 344.8000 ;
      RECT 209.0500 344.1000 209.5500 344.8000 ;
      RECT 208.2500 344.1000 208.7500 344.8000 ;
      RECT 207.4500 344.1000 207.9500 344.8000 ;
      RECT 206.6500 344.1000 207.1500 344.8000 ;
      RECT 205.8500 344.1000 206.3500 344.8000 ;
      RECT 205.0500 344.1000 205.5500 344.8000 ;
      RECT 204.2500 344.1000 204.7500 344.8000 ;
      RECT 203.4500 344.1000 203.9500 344.8000 ;
      RECT 202.6500 344.1000 203.1500 344.8000 ;
      RECT 201.8500 344.1000 202.3500 344.8000 ;
      RECT 201.0500 344.1000 201.5500 344.8000 ;
      RECT 200.2500 344.1000 200.7500 344.8000 ;
      RECT 199.4500 344.1000 199.9500 344.8000 ;
      RECT 198.6500 344.1000 199.1500 344.8000 ;
      RECT 197.8500 344.1000 198.3500 344.8000 ;
      RECT 197.0500 344.1000 197.5500 344.8000 ;
      RECT 196.2500 344.1000 196.7500 344.8000 ;
      RECT 195.4500 344.1000 195.9500 344.8000 ;
      RECT 194.6500 344.1000 195.1500 344.8000 ;
      RECT 193.8500 344.1000 194.3500 344.8000 ;
      RECT 193.0500 344.1000 193.5500 344.8000 ;
      RECT 192.2500 344.1000 192.7500 344.8000 ;
      RECT 191.4500 344.1000 191.9500 344.8000 ;
      RECT 190.6500 344.1000 191.1500 344.8000 ;
      RECT 189.8500 344.1000 190.3500 344.8000 ;
      RECT 189.0500 344.1000 189.5500 344.8000 ;
      RECT 188.2500 344.1000 188.7500 344.8000 ;
      RECT 187.4500 344.1000 187.9500 344.8000 ;
      RECT 186.6500 344.1000 187.1500 344.8000 ;
      RECT 185.8500 344.1000 186.3500 344.8000 ;
      RECT 185.0500 344.1000 185.5500 344.8000 ;
      RECT 184.2500 344.1000 184.7500 344.8000 ;
      RECT 183.4500 344.1000 183.9500 344.8000 ;
      RECT 182.6500 344.1000 183.1500 344.8000 ;
      RECT 181.8500 344.1000 182.3500 344.8000 ;
      RECT 181.0500 344.1000 181.5500 344.8000 ;
      RECT 180.2500 344.1000 180.7500 344.8000 ;
      RECT 179.4500 344.1000 179.9500 344.8000 ;
      RECT 178.6500 344.1000 179.1500 344.8000 ;
      RECT 177.8500 344.1000 178.3500 344.8000 ;
      RECT 177.0500 344.1000 177.5500 344.8000 ;
      RECT 176.2500 344.1000 176.7500 344.8000 ;
      RECT 175.4500 344.1000 175.9500 344.8000 ;
      RECT 174.6500 344.1000 175.1500 344.8000 ;
      RECT 173.8500 344.1000 174.3500 344.8000 ;
      RECT 173.0500 344.1000 173.5500 344.8000 ;
      RECT 172.2500 344.1000 172.7500 344.8000 ;
      RECT 171.4500 344.1000 171.9500 344.8000 ;
      RECT 170.6500 344.1000 171.1500 344.8000 ;
      RECT 169.8500 344.1000 170.3500 344.8000 ;
      RECT 169.0500 344.1000 169.5500 344.8000 ;
      RECT 168.2500 344.1000 168.7500 344.8000 ;
      RECT 167.4500 344.1000 167.9500 344.8000 ;
      RECT 166.6500 344.1000 167.1500 344.8000 ;
      RECT 165.8500 344.1000 166.3500 344.8000 ;
      RECT 165.0500 344.1000 165.5500 344.8000 ;
      RECT 164.2500 344.1000 164.7500 344.8000 ;
      RECT 163.4500 344.1000 163.9500 344.8000 ;
      RECT 162.6500 344.1000 163.1500 344.8000 ;
      RECT 161.8500 344.1000 162.3500 344.8000 ;
      RECT 161.0500 344.1000 161.5500 344.8000 ;
      RECT 160.2500 344.1000 160.7500 344.8000 ;
      RECT 159.4500 344.1000 159.9500 344.8000 ;
      RECT 158.6500 344.1000 159.1500 344.8000 ;
      RECT 157.8500 344.1000 158.3500 344.8000 ;
      RECT 157.0500 344.1000 157.5500 344.8000 ;
      RECT 156.2500 344.1000 156.7500 344.8000 ;
      RECT 155.4500 344.1000 155.9500 344.8000 ;
      RECT 154.6500 344.1000 155.1500 344.8000 ;
      RECT 153.8500 344.1000 154.3500 344.8000 ;
      RECT 153.0500 344.1000 153.5500 344.8000 ;
      RECT 152.2500 344.1000 152.7500 344.8000 ;
      RECT 151.4500 344.1000 151.9500 344.8000 ;
      RECT 150.6500 344.1000 151.1500 344.8000 ;
      RECT 149.8500 344.1000 150.3500 344.8000 ;
      RECT 149.0500 344.1000 149.5500 344.8000 ;
      RECT 148.2500 344.1000 148.7500 344.8000 ;
      RECT 147.4500 344.1000 147.9500 344.8000 ;
      RECT 146.6500 344.1000 147.1500 344.8000 ;
      RECT 145.8500 344.1000 146.3500 344.8000 ;
      RECT 145.0500 344.1000 145.5500 344.8000 ;
      RECT 144.2500 344.1000 144.7500 344.8000 ;
      RECT 143.4500 344.1000 143.9500 344.8000 ;
      RECT 142.6500 344.1000 143.1500 344.8000 ;
      RECT 141.8500 344.1000 142.3500 344.8000 ;
      RECT 141.0500 344.1000 141.5500 344.8000 ;
      RECT 140.2500 344.1000 140.7500 344.8000 ;
      RECT 139.4500 344.1000 139.9500 344.8000 ;
      RECT 138.6500 344.1000 139.1500 344.8000 ;
      RECT 137.8500 344.1000 138.3500 344.8000 ;
      RECT 137.0500 344.1000 137.5500 344.8000 ;
      RECT 136.2500 344.1000 136.7500 344.8000 ;
      RECT 135.4500 344.1000 135.9500 344.8000 ;
      RECT 134.6500 344.1000 135.1500 344.8000 ;
      RECT 133.8500 344.1000 134.3500 344.8000 ;
      RECT 133.0500 344.1000 133.5500 344.8000 ;
      RECT 132.2500 344.1000 132.7500 344.8000 ;
      RECT 131.4500 344.1000 131.9500 344.8000 ;
      RECT 130.6500 344.1000 131.1500 344.8000 ;
      RECT 129.8500 344.1000 130.3500 344.8000 ;
      RECT 129.0500 344.1000 129.5500 344.8000 ;
      RECT 128.2500 344.1000 128.7500 344.8000 ;
      RECT 127.4500 344.1000 127.9500 344.8000 ;
      RECT 126.6500 344.1000 127.1500 344.8000 ;
      RECT 125.8500 344.1000 126.3500 344.8000 ;
      RECT 125.0500 344.1000 125.5500 344.8000 ;
      RECT 124.2500 344.1000 124.7500 344.8000 ;
      RECT 123.4500 344.1000 123.9500 344.8000 ;
      RECT 122.6500 344.1000 123.1500 344.8000 ;
      RECT 0.0000 344.1000 122.3500 344.8000 ;
      RECT 0.0000 0.7000 346.4000 344.1000 ;
      RECT 224.2500 0.0000 346.4000 0.7000 ;
      RECT 223.4500 0.0000 223.9500 0.7000 ;
      RECT 222.6500 0.0000 223.1500 0.7000 ;
      RECT 221.8500 0.0000 222.3500 0.7000 ;
      RECT 221.0500 0.0000 221.5500 0.7000 ;
      RECT 220.2500 0.0000 220.7500 0.7000 ;
      RECT 219.4500 0.0000 219.9500 0.7000 ;
      RECT 218.6500 0.0000 219.1500 0.7000 ;
      RECT 217.8500 0.0000 218.3500 0.7000 ;
      RECT 217.0500 0.0000 217.5500 0.7000 ;
      RECT 216.2500 0.0000 216.7500 0.7000 ;
      RECT 215.4500 0.0000 215.9500 0.7000 ;
      RECT 214.6500 0.0000 215.1500 0.7000 ;
      RECT 213.8500 0.0000 214.3500 0.7000 ;
      RECT 213.0500 0.0000 213.5500 0.7000 ;
      RECT 212.2500 0.0000 212.7500 0.7000 ;
      RECT 211.4500 0.0000 211.9500 0.7000 ;
      RECT 210.6500 0.0000 211.1500 0.7000 ;
      RECT 209.8500 0.0000 210.3500 0.7000 ;
      RECT 209.0500 0.0000 209.5500 0.7000 ;
      RECT 208.2500 0.0000 208.7500 0.7000 ;
      RECT 207.4500 0.0000 207.9500 0.7000 ;
      RECT 206.6500 0.0000 207.1500 0.7000 ;
      RECT 205.8500 0.0000 206.3500 0.7000 ;
      RECT 205.0500 0.0000 205.5500 0.7000 ;
      RECT 204.2500 0.0000 204.7500 0.7000 ;
      RECT 203.4500 0.0000 203.9500 0.7000 ;
      RECT 202.6500 0.0000 203.1500 0.7000 ;
      RECT 201.8500 0.0000 202.3500 0.7000 ;
      RECT 201.0500 0.0000 201.5500 0.7000 ;
      RECT 200.2500 0.0000 200.7500 0.7000 ;
      RECT 199.4500 0.0000 199.9500 0.7000 ;
      RECT 198.6500 0.0000 199.1500 0.7000 ;
      RECT 197.8500 0.0000 198.3500 0.7000 ;
      RECT 197.0500 0.0000 197.5500 0.7000 ;
      RECT 196.2500 0.0000 196.7500 0.7000 ;
      RECT 195.4500 0.0000 195.9500 0.7000 ;
      RECT 194.6500 0.0000 195.1500 0.7000 ;
      RECT 193.8500 0.0000 194.3500 0.7000 ;
      RECT 193.0500 0.0000 193.5500 0.7000 ;
      RECT 192.2500 0.0000 192.7500 0.7000 ;
      RECT 191.4500 0.0000 191.9500 0.7000 ;
      RECT 190.6500 0.0000 191.1500 0.7000 ;
      RECT 189.8500 0.0000 190.3500 0.7000 ;
      RECT 189.0500 0.0000 189.5500 0.7000 ;
      RECT 188.2500 0.0000 188.7500 0.7000 ;
      RECT 187.4500 0.0000 187.9500 0.7000 ;
      RECT 186.6500 0.0000 187.1500 0.7000 ;
      RECT 185.8500 0.0000 186.3500 0.7000 ;
      RECT 185.0500 0.0000 185.5500 0.7000 ;
      RECT 184.2500 0.0000 184.7500 0.7000 ;
      RECT 183.4500 0.0000 183.9500 0.7000 ;
      RECT 182.6500 0.0000 183.1500 0.7000 ;
      RECT 181.8500 0.0000 182.3500 0.7000 ;
      RECT 181.0500 0.0000 181.5500 0.7000 ;
      RECT 180.2500 0.0000 180.7500 0.7000 ;
      RECT 179.4500 0.0000 179.9500 0.7000 ;
      RECT 178.6500 0.0000 179.1500 0.7000 ;
      RECT 177.8500 0.0000 178.3500 0.7000 ;
      RECT 177.0500 0.0000 177.5500 0.7000 ;
      RECT 176.2500 0.0000 176.7500 0.7000 ;
      RECT 175.4500 0.0000 175.9500 0.7000 ;
      RECT 174.6500 0.0000 175.1500 0.7000 ;
      RECT 173.8500 0.0000 174.3500 0.7000 ;
      RECT 173.0500 0.0000 173.5500 0.7000 ;
      RECT 172.2500 0.0000 172.7500 0.7000 ;
      RECT 171.4500 0.0000 171.9500 0.7000 ;
      RECT 170.6500 0.0000 171.1500 0.7000 ;
      RECT 169.8500 0.0000 170.3500 0.7000 ;
      RECT 169.0500 0.0000 169.5500 0.7000 ;
      RECT 168.2500 0.0000 168.7500 0.7000 ;
      RECT 167.4500 0.0000 167.9500 0.7000 ;
      RECT 166.6500 0.0000 167.1500 0.7000 ;
      RECT 165.8500 0.0000 166.3500 0.7000 ;
      RECT 165.0500 0.0000 165.5500 0.7000 ;
      RECT 164.2500 0.0000 164.7500 0.7000 ;
      RECT 163.4500 0.0000 163.9500 0.7000 ;
      RECT 162.6500 0.0000 163.1500 0.7000 ;
      RECT 161.8500 0.0000 162.3500 0.7000 ;
      RECT 161.0500 0.0000 161.5500 0.7000 ;
      RECT 160.2500 0.0000 160.7500 0.7000 ;
      RECT 159.4500 0.0000 159.9500 0.7000 ;
      RECT 158.6500 0.0000 159.1500 0.7000 ;
      RECT 157.8500 0.0000 158.3500 0.7000 ;
      RECT 157.0500 0.0000 157.5500 0.7000 ;
      RECT 156.2500 0.0000 156.7500 0.7000 ;
      RECT 155.4500 0.0000 155.9500 0.7000 ;
      RECT 154.6500 0.0000 155.1500 0.7000 ;
      RECT 153.8500 0.0000 154.3500 0.7000 ;
      RECT 153.0500 0.0000 153.5500 0.7000 ;
      RECT 152.2500 0.0000 152.7500 0.7000 ;
      RECT 151.4500 0.0000 151.9500 0.7000 ;
      RECT 150.6500 0.0000 151.1500 0.7000 ;
      RECT 149.8500 0.0000 150.3500 0.7000 ;
      RECT 149.0500 0.0000 149.5500 0.7000 ;
      RECT 148.2500 0.0000 148.7500 0.7000 ;
      RECT 147.4500 0.0000 147.9500 0.7000 ;
      RECT 146.6500 0.0000 147.1500 0.7000 ;
      RECT 145.8500 0.0000 146.3500 0.7000 ;
      RECT 145.0500 0.0000 145.5500 0.7000 ;
      RECT 144.2500 0.0000 144.7500 0.7000 ;
      RECT 143.4500 0.0000 143.9500 0.7000 ;
      RECT 142.6500 0.0000 143.1500 0.7000 ;
      RECT 141.8500 0.0000 142.3500 0.7000 ;
      RECT 141.0500 0.0000 141.5500 0.7000 ;
      RECT 140.2500 0.0000 140.7500 0.7000 ;
      RECT 139.4500 0.0000 139.9500 0.7000 ;
      RECT 138.6500 0.0000 139.1500 0.7000 ;
      RECT 137.8500 0.0000 138.3500 0.7000 ;
      RECT 137.0500 0.0000 137.5500 0.7000 ;
      RECT 136.2500 0.0000 136.7500 0.7000 ;
      RECT 135.4500 0.0000 135.9500 0.7000 ;
      RECT 134.6500 0.0000 135.1500 0.7000 ;
      RECT 133.8500 0.0000 134.3500 0.7000 ;
      RECT 133.0500 0.0000 133.5500 0.7000 ;
      RECT 132.2500 0.0000 132.7500 0.7000 ;
      RECT 131.4500 0.0000 131.9500 0.7000 ;
      RECT 130.6500 0.0000 131.1500 0.7000 ;
      RECT 129.8500 0.0000 130.3500 0.7000 ;
      RECT 129.0500 0.0000 129.5500 0.7000 ;
      RECT 128.2500 0.0000 128.7500 0.7000 ;
      RECT 127.4500 0.0000 127.9500 0.7000 ;
      RECT 126.6500 0.0000 127.1500 0.7000 ;
      RECT 125.8500 0.0000 126.3500 0.7000 ;
      RECT 125.0500 0.0000 125.5500 0.7000 ;
      RECT 124.2500 0.0000 124.7500 0.7000 ;
      RECT 123.4500 0.0000 123.9500 0.7000 ;
      RECT 122.6500 0.0000 123.1500 0.7000 ;
      RECT 0.0000 0.0000 122.3500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 20.9500 346.4000 344.8000 ;
      RECT 0.7000 20.6500 346.4000 20.9500 ;
      RECT 0.0000 20.1500 346.4000 20.6500 ;
      RECT 0.7000 19.8500 346.4000 20.1500 ;
      RECT 0.0000 19.3500 346.4000 19.8500 ;
      RECT 0.7000 19.0500 346.4000 19.3500 ;
      RECT 0.0000 18.5500 346.4000 19.0500 ;
      RECT 0.7000 18.2500 346.4000 18.5500 ;
      RECT 0.0000 17.7500 346.4000 18.2500 ;
      RECT 0.7000 17.4500 346.4000 17.7500 ;
      RECT 0.0000 16.9500 346.4000 17.4500 ;
      RECT 0.7000 16.6500 346.4000 16.9500 ;
      RECT 0.0000 16.1500 346.4000 16.6500 ;
      RECT 0.7000 15.8500 346.4000 16.1500 ;
      RECT 0.0000 0.0000 346.4000 15.8500 ;
    LAYER M4 ;
      RECT 0.0000 295.4650 346.4000 344.8000 ;
      RECT 288.8850 295.3000 346.4000 295.4650 ;
      RECT 262.6200 295.3000 285.8850 295.4650 ;
      RECT 236.3550 295.3000 259.6200 295.4650 ;
      RECT 210.0900 295.3000 233.3550 295.4650 ;
      RECT 183.8250 295.3000 207.0900 295.4650 ;
      RECT 157.5600 295.3000 180.8250 295.4650 ;
      RECT 131.2950 295.3000 154.5600 295.4650 ;
      RECT 105.0300 295.3000 128.2950 295.4650 ;
      RECT 78.7650 295.3000 102.0300 295.4650 ;
      RECT 52.5000 295.3000 75.7650 295.4650 ;
      RECT 296.8850 49.5000 346.4000 295.3000 ;
      RECT 288.8850 49.5000 293.8850 295.3000 ;
      RECT 270.6200 49.5000 285.8850 295.3000 ;
      RECT 262.6200 49.5000 267.6200 295.3000 ;
      RECT 244.3550 49.5000 259.6200 295.3000 ;
      RECT 236.3550 49.5000 241.3550 295.3000 ;
      RECT 218.0900 49.5000 233.3550 295.3000 ;
      RECT 210.0900 49.5000 215.0900 295.3000 ;
      RECT 191.8250 49.5000 207.0900 295.3000 ;
      RECT 183.8250 49.5000 188.8250 295.3000 ;
      RECT 165.5600 49.5000 180.8250 295.3000 ;
      RECT 157.5600 49.5000 162.5600 295.3000 ;
      RECT 139.2950 49.5000 154.5600 295.3000 ;
      RECT 131.2950 49.5000 136.2950 295.3000 ;
      RECT 113.0300 49.5000 128.2950 295.3000 ;
      RECT 105.0300 49.5000 110.0300 295.3000 ;
      RECT 86.7650 49.5000 102.0300 295.3000 ;
      RECT 78.7650 49.5000 83.7650 295.3000 ;
      RECT 60.5000 49.5000 75.7650 295.3000 ;
      RECT 52.5000 49.5000 57.5000 295.3000 ;
      RECT 288.8850 49.3350 346.4000 49.5000 ;
      RECT 262.6200 49.3350 285.8850 49.5000 ;
      RECT 236.3550 49.3350 259.6200 49.5000 ;
      RECT 210.0900 49.3350 233.3550 49.5000 ;
      RECT 183.8250 49.3350 207.0900 49.5000 ;
      RECT 157.5600 49.3350 180.8250 49.5000 ;
      RECT 131.2950 49.3350 154.5600 49.5000 ;
      RECT 105.0300 49.3350 128.2950 49.5000 ;
      RECT 78.7650 49.3350 102.0300 49.5000 ;
      RECT 52.5000 49.3350 75.7650 49.5000 ;
      RECT 0.0000 49.3350 49.5000 295.4650 ;
      RECT 0.0000 0.0000 346.4000 49.3350 ;
  END
END sram_w16

END LIBRARY
