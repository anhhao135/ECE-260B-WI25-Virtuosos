##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Mon Mar 10 10:44:14 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO mac_8in
  CLASS BLOCK ;
  SIZE 160.6000 BY 158.6000 ;
  FOREIGN mac_8in 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 90.4500 0.0000 90.5500 0.6000 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 89.4500 0.0000 89.5500 0.6000 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 88.4500 0.0000 88.5500 0.6000 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 87.4500 0.0000 87.5500 0.6000 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 86.4500 0.0000 86.5500 0.6000 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 85.4500 0.0000 85.5500 0.6000 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 84.4500 0.0000 84.5500 0.6000 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 83.4500 0.0000 83.5500 0.6000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 82.4500 0.0000 82.5500 0.6000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 81.4500 0.0000 81.5500 0.6000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 80.4500 0.0000 80.5500 0.6000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 79.4500 0.0000 79.5500 0.6000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 78.4500 0.0000 78.5500 0.6000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 77.4500 0.0000 77.5500 0.6000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 76.4500 0.0000 76.5500 0.6000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 75.4500 0.0000 75.5500 0.6000 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 74.4500 0.0000 74.5500 0.6000 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 73.4500 0.0000 73.5500 0.6000 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 72.4500 0.0000 72.5500 0.6000 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 71.4500 0.0000 71.5500 0.6000 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 70.4500 0.0000 70.5500 0.6000 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 69.4500 0.0000 69.5500 0.6000 ;
    END
  END out[0]
  PIN a[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 77.5500 0.6000 77.6500 ;
    END
  END a[63]
  PIN a[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 76.5500 0.6000 76.6500 ;
    END
  END a[62]
  PIN a[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 75.5500 0.6000 75.6500 ;
    END
  END a[61]
  PIN a[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 74.5500 0.6000 74.6500 ;
    END
  END a[60]
  PIN a[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 73.5500 0.6000 73.6500 ;
    END
  END a[59]
  PIN a[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.5500 0.6000 72.6500 ;
    END
  END a[58]
  PIN a[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 71.5500 0.6000 71.6500 ;
    END
  END a[57]
  PIN a[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 70.5500 0.6000 70.6500 ;
    END
  END a[56]
  PIN a[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.5500 0.6000 69.6500 ;
    END
  END a[55]
  PIN a[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 68.5500 0.6000 68.6500 ;
    END
  END a[54]
  PIN a[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 67.5500 0.6000 67.6500 ;
    END
  END a[53]
  PIN a[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 66.5500 0.6000 66.6500 ;
    END
  END a[52]
  PIN a[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.5500 0.6000 65.6500 ;
    END
  END a[51]
  PIN a[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.5500 0.6000 64.6500 ;
    END
  END a[50]
  PIN a[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.5500 0.6000 63.6500 ;
    END
  END a[49]
  PIN a[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.5500 0.6000 62.6500 ;
    END
  END a[48]
  PIN a[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.5500 0.6000 61.6500 ;
    END
  END a[47]
  PIN a[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.5500 0.6000 60.6500 ;
    END
  END a[46]
  PIN a[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.5500 0.6000 59.6500 ;
    END
  END a[45]
  PIN a[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 58.5500 0.6000 58.6500 ;
    END
  END a[44]
  PIN a[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.5500 0.6000 57.6500 ;
    END
  END a[43]
  PIN a[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.5500 0.6000 56.6500 ;
    END
  END a[42]
  PIN a[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.5500 0.6000 55.6500 ;
    END
  END a[41]
  PIN a[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.5500 0.6000 54.6500 ;
    END
  END a[40]
  PIN a[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.5500 0.6000 53.6500 ;
    END
  END a[39]
  PIN a[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.5500 0.6000 52.6500 ;
    END
  END a[38]
  PIN a[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.5500 0.6000 51.6500 ;
    END
  END a[37]
  PIN a[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 50.5500 0.6000 50.6500 ;
    END
  END a[36]
  PIN a[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.5500 0.6000 49.6500 ;
    END
  END a[35]
  PIN a[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.5500 0.6000 48.6500 ;
    END
  END a[34]
  PIN a[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 47.5500 0.6000 47.6500 ;
    END
  END a[33]
  PIN a[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 46.5500 0.6000 46.6500 ;
    END
  END a[32]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 45.5500 0.6000 45.6500 ;
    END
  END a[31]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 44.5500 0.6000 44.6500 ;
    END
  END a[30]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 43.5500 0.6000 43.6500 ;
    END
  END a[29]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 42.5500 0.6000 42.6500 ;
    END
  END a[28]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 41.5500 0.6000 41.6500 ;
    END
  END a[27]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 40.5500 0.6000 40.6500 ;
    END
  END a[26]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 39.5500 0.6000 39.6500 ;
    END
  END a[25]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 38.5500 0.6000 38.6500 ;
    END
  END a[24]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 37.5500 0.6000 37.6500 ;
    END
  END a[23]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 36.5500 0.6000 36.6500 ;
    END
  END a[22]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 35.5500 0.6000 35.6500 ;
    END
  END a[21]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.5500 0.6000 34.6500 ;
    END
  END a[20]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 33.5500 0.6000 33.6500 ;
    END
  END a[19]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 32.5500 0.6000 32.6500 ;
    END
  END a[18]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 31.5500 0.6000 31.6500 ;
    END
  END a[17]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 30.5500 0.6000 30.6500 ;
    END
  END a[16]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 29.5500 0.6000 29.6500 ;
    END
  END a[15]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 28.5500 0.6000 28.6500 ;
    END
  END a[14]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 27.5500 0.6000 27.6500 ;
    END
  END a[13]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 26.5500 0.6000 26.6500 ;
    END
  END a[12]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 25.5500 0.6000 25.6500 ;
    END
  END a[11]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 24.5500 0.6000 24.6500 ;
    END
  END a[10]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 23.5500 0.6000 23.6500 ;
    END
  END a[9]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 22.5500 0.6000 22.6500 ;
    END
  END a[8]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 21.5500 0.6000 21.6500 ;
    END
  END a[7]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.5500 0.6000 20.6500 ;
    END
  END a[6]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.5500 0.6000 19.6500 ;
    END
  END a[5]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.5500 0.6000 18.6500 ;
    END
  END a[4]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.5500 0.6000 17.6500 ;
    END
  END a[3]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.5500 0.6000 16.6500 ;
    END
  END a[2]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.5500 0.6000 15.6500 ;
    END
  END a[1]
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 14.5500 0.6000 14.6500 ;
    END
  END a[0]
  PIN b[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 141.5500 0.6000 141.6500 ;
    END
  END b[63]
  PIN b[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 140.5500 0.6000 140.6500 ;
    END
  END b[62]
  PIN b[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 139.5500 0.6000 139.6500 ;
    END
  END b[61]
  PIN b[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 138.5500 0.6000 138.6500 ;
    END
  END b[60]
  PIN b[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 137.5500 0.6000 137.6500 ;
    END
  END b[59]
  PIN b[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 136.5500 0.6000 136.6500 ;
    END
  END b[58]
  PIN b[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 135.5500 0.6000 135.6500 ;
    END
  END b[57]
  PIN b[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 134.5500 0.6000 134.6500 ;
    END
  END b[56]
  PIN b[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 133.5500 0.6000 133.6500 ;
    END
  END b[55]
  PIN b[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 132.5500 0.6000 132.6500 ;
    END
  END b[54]
  PIN b[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 131.5500 0.6000 131.6500 ;
    END
  END b[53]
  PIN b[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 130.5500 0.6000 130.6500 ;
    END
  END b[52]
  PIN b[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 129.5500 0.6000 129.6500 ;
    END
  END b[51]
  PIN b[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 128.5500 0.6000 128.6500 ;
    END
  END b[50]
  PIN b[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 127.5500 0.6000 127.6500 ;
    END
  END b[49]
  PIN b[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 126.5500 0.6000 126.6500 ;
    END
  END b[48]
  PIN b[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 125.5500 0.6000 125.6500 ;
    END
  END b[47]
  PIN b[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 124.5500 0.6000 124.6500 ;
    END
  END b[46]
  PIN b[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 123.5500 0.6000 123.6500 ;
    END
  END b[45]
  PIN b[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 122.5500 0.6000 122.6500 ;
    END
  END b[44]
  PIN b[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 121.5500 0.6000 121.6500 ;
    END
  END b[43]
  PIN b[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 120.5500 0.6000 120.6500 ;
    END
  END b[42]
  PIN b[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 119.5500 0.6000 119.6500 ;
    END
  END b[41]
  PIN b[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 118.5500 0.6000 118.6500 ;
    END
  END b[40]
  PIN b[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 117.5500 0.6000 117.6500 ;
    END
  END b[39]
  PIN b[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 116.5500 0.6000 116.6500 ;
    END
  END b[38]
  PIN b[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 115.5500 0.6000 115.6500 ;
    END
  END b[37]
  PIN b[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 114.5500 0.6000 114.6500 ;
    END
  END b[36]
  PIN b[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 113.5500 0.6000 113.6500 ;
    END
  END b[35]
  PIN b[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 112.5500 0.6000 112.6500 ;
    END
  END b[34]
  PIN b[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 111.5500 0.6000 111.6500 ;
    END
  END b[33]
  PIN b[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 110.5500 0.6000 110.6500 ;
    END
  END b[32]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 109.5500 0.6000 109.6500 ;
    END
  END b[31]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 108.5500 0.6000 108.6500 ;
    END
  END b[30]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 107.5500 0.6000 107.6500 ;
    END
  END b[29]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 106.5500 0.6000 106.6500 ;
    END
  END b[28]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 105.5500 0.6000 105.6500 ;
    END
  END b[27]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 104.5500 0.6000 104.6500 ;
    END
  END b[26]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 103.5500 0.6000 103.6500 ;
    END
  END b[25]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 102.5500 0.6000 102.6500 ;
    END
  END b[24]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 101.5500 0.6000 101.6500 ;
    END
  END b[23]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 100.5500 0.6000 100.6500 ;
    END
  END b[22]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 99.5500 0.6000 99.6500 ;
    END
  END b[21]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 98.5500 0.6000 98.6500 ;
    END
  END b[20]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 97.5500 0.6000 97.6500 ;
    END
  END b[19]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.5500 0.6000 96.6500 ;
    END
  END b[18]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 95.5500 0.6000 95.6500 ;
    END
  END b[17]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 94.5500 0.6000 94.6500 ;
    END
  END b[16]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 93.5500 0.6000 93.6500 ;
    END
  END b[15]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 92.5500 0.6000 92.6500 ;
    END
  END b[14]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 91.5500 0.6000 91.6500 ;
    END
  END b[13]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 90.5500 0.6000 90.6500 ;
    END
  END b[12]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 89.5500 0.6000 89.6500 ;
    END
  END b[11]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 88.5500 0.6000 88.6500 ;
    END
  END b[10]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 87.5500 0.6000 87.6500 ;
    END
  END b[9]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 86.5500 0.6000 86.6500 ;
    END
  END b[8]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 85.5500 0.6000 85.6500 ;
    END
  END b[7]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 84.5500 0.6000 84.6500 ;
    END
  END b[6]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 83.5500 0.6000 83.6500 ;
    END
  END b[5]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 82.5500 0.6000 82.6500 ;
    END
  END b[4]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 81.5500 0.6000 81.6500 ;
    END
  END b[3]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 80.5500 0.6000 80.6500 ;
    END
  END b[2]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 79.5500 0.6000 79.6500 ;
    END
  END b[1]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 78.5500 0.6000 78.6500 ;
    END
  END b[0]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 142.5500 0.6000 142.6500 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 143.5500 0.6000 143.6500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M3 ;
      RECT 0.0000 143.7500 160.6000 158.6000 ;
      RECT 0.7000 143.4500 160.6000 143.7500 ;
      RECT 0.0000 142.7500 160.6000 143.4500 ;
      RECT 0.7000 142.4500 160.6000 142.7500 ;
      RECT 0.0000 141.7500 160.6000 142.4500 ;
      RECT 0.7000 141.4500 160.6000 141.7500 ;
      RECT 0.0000 140.7500 160.6000 141.4500 ;
      RECT 0.7000 140.4500 160.6000 140.7500 ;
      RECT 0.0000 139.7500 160.6000 140.4500 ;
      RECT 0.7000 139.4500 160.6000 139.7500 ;
      RECT 0.0000 138.7500 160.6000 139.4500 ;
      RECT 0.7000 138.4500 160.6000 138.7500 ;
      RECT 0.0000 137.7500 160.6000 138.4500 ;
      RECT 0.7000 137.4500 160.6000 137.7500 ;
      RECT 0.0000 136.7500 160.6000 137.4500 ;
      RECT 0.7000 136.4500 160.6000 136.7500 ;
      RECT 0.0000 135.7500 160.6000 136.4500 ;
      RECT 0.7000 135.4500 160.6000 135.7500 ;
      RECT 0.0000 134.7500 160.6000 135.4500 ;
      RECT 0.7000 134.4500 160.6000 134.7500 ;
      RECT 0.0000 133.7500 160.6000 134.4500 ;
      RECT 0.7000 133.4500 160.6000 133.7500 ;
      RECT 0.0000 132.7500 160.6000 133.4500 ;
      RECT 0.7000 132.4500 160.6000 132.7500 ;
      RECT 0.0000 131.7500 160.6000 132.4500 ;
      RECT 0.7000 131.4500 160.6000 131.7500 ;
      RECT 0.0000 130.7500 160.6000 131.4500 ;
      RECT 0.7000 130.4500 160.6000 130.7500 ;
      RECT 0.0000 129.7500 160.6000 130.4500 ;
      RECT 0.7000 129.4500 160.6000 129.7500 ;
      RECT 0.0000 128.7500 160.6000 129.4500 ;
      RECT 0.7000 128.4500 160.6000 128.7500 ;
      RECT 0.0000 127.7500 160.6000 128.4500 ;
      RECT 0.7000 127.4500 160.6000 127.7500 ;
      RECT 0.0000 126.7500 160.6000 127.4500 ;
      RECT 0.7000 126.4500 160.6000 126.7500 ;
      RECT 0.0000 125.7500 160.6000 126.4500 ;
      RECT 0.7000 125.4500 160.6000 125.7500 ;
      RECT 0.0000 124.7500 160.6000 125.4500 ;
      RECT 0.7000 124.4500 160.6000 124.7500 ;
      RECT 0.0000 123.7500 160.6000 124.4500 ;
      RECT 0.7000 123.4500 160.6000 123.7500 ;
      RECT 0.0000 122.7500 160.6000 123.4500 ;
      RECT 0.7000 122.4500 160.6000 122.7500 ;
      RECT 0.0000 121.7500 160.6000 122.4500 ;
      RECT 0.7000 121.4500 160.6000 121.7500 ;
      RECT 0.0000 120.7500 160.6000 121.4500 ;
      RECT 0.7000 120.4500 160.6000 120.7500 ;
      RECT 0.0000 119.7500 160.6000 120.4500 ;
      RECT 0.7000 119.4500 160.6000 119.7500 ;
      RECT 0.0000 118.7500 160.6000 119.4500 ;
      RECT 0.7000 118.4500 160.6000 118.7500 ;
      RECT 0.0000 117.7500 160.6000 118.4500 ;
      RECT 0.7000 117.4500 160.6000 117.7500 ;
      RECT 0.0000 116.7500 160.6000 117.4500 ;
      RECT 0.7000 116.4500 160.6000 116.7500 ;
      RECT 0.0000 115.7500 160.6000 116.4500 ;
      RECT 0.7000 115.4500 160.6000 115.7500 ;
      RECT 0.0000 114.7500 160.6000 115.4500 ;
      RECT 0.7000 114.4500 160.6000 114.7500 ;
      RECT 0.0000 113.7500 160.6000 114.4500 ;
      RECT 0.7000 113.4500 160.6000 113.7500 ;
      RECT 0.0000 112.7500 160.6000 113.4500 ;
      RECT 0.7000 112.4500 160.6000 112.7500 ;
      RECT 0.0000 111.7500 160.6000 112.4500 ;
      RECT 0.7000 111.4500 160.6000 111.7500 ;
      RECT 0.0000 110.7500 160.6000 111.4500 ;
      RECT 0.7000 110.4500 160.6000 110.7500 ;
      RECT 0.0000 109.7500 160.6000 110.4500 ;
      RECT 0.7000 109.4500 160.6000 109.7500 ;
      RECT 0.0000 108.7500 160.6000 109.4500 ;
      RECT 0.7000 108.4500 160.6000 108.7500 ;
      RECT 0.0000 107.7500 160.6000 108.4500 ;
      RECT 0.7000 107.4500 160.6000 107.7500 ;
      RECT 0.0000 106.7500 160.6000 107.4500 ;
      RECT 0.7000 106.4500 160.6000 106.7500 ;
      RECT 0.0000 105.7500 160.6000 106.4500 ;
      RECT 0.7000 105.4500 160.6000 105.7500 ;
      RECT 0.0000 104.7500 160.6000 105.4500 ;
      RECT 0.7000 104.4500 160.6000 104.7500 ;
      RECT 0.0000 103.7500 160.6000 104.4500 ;
      RECT 0.7000 103.4500 160.6000 103.7500 ;
      RECT 0.0000 102.7500 160.6000 103.4500 ;
      RECT 0.7000 102.4500 160.6000 102.7500 ;
      RECT 0.0000 101.7500 160.6000 102.4500 ;
      RECT 0.7000 101.4500 160.6000 101.7500 ;
      RECT 0.0000 100.7500 160.6000 101.4500 ;
      RECT 0.7000 100.4500 160.6000 100.7500 ;
      RECT 0.0000 99.7500 160.6000 100.4500 ;
      RECT 0.7000 99.4500 160.6000 99.7500 ;
      RECT 0.0000 98.7500 160.6000 99.4500 ;
      RECT 0.7000 98.4500 160.6000 98.7500 ;
      RECT 0.0000 97.7500 160.6000 98.4500 ;
      RECT 0.7000 97.4500 160.6000 97.7500 ;
      RECT 0.0000 96.7500 160.6000 97.4500 ;
      RECT 0.7000 96.4500 160.6000 96.7500 ;
      RECT 0.0000 95.7500 160.6000 96.4500 ;
      RECT 0.7000 95.4500 160.6000 95.7500 ;
      RECT 0.0000 94.7500 160.6000 95.4500 ;
      RECT 0.7000 94.4500 160.6000 94.7500 ;
      RECT 0.0000 93.7500 160.6000 94.4500 ;
      RECT 0.7000 93.4500 160.6000 93.7500 ;
      RECT 0.0000 92.7500 160.6000 93.4500 ;
      RECT 0.7000 92.4500 160.6000 92.7500 ;
      RECT 0.0000 91.7500 160.6000 92.4500 ;
      RECT 0.7000 91.4500 160.6000 91.7500 ;
      RECT 0.0000 90.7500 160.6000 91.4500 ;
      RECT 0.7000 90.4500 160.6000 90.7500 ;
      RECT 0.0000 89.7500 160.6000 90.4500 ;
      RECT 0.7000 89.4500 160.6000 89.7500 ;
      RECT 0.0000 88.7500 160.6000 89.4500 ;
      RECT 0.7000 88.4500 160.6000 88.7500 ;
      RECT 0.0000 87.7500 160.6000 88.4500 ;
      RECT 0.7000 87.4500 160.6000 87.7500 ;
      RECT 0.0000 86.7500 160.6000 87.4500 ;
      RECT 0.7000 86.4500 160.6000 86.7500 ;
      RECT 0.0000 85.7500 160.6000 86.4500 ;
      RECT 0.7000 85.4500 160.6000 85.7500 ;
      RECT 0.0000 84.7500 160.6000 85.4500 ;
      RECT 0.7000 84.4500 160.6000 84.7500 ;
      RECT 0.0000 83.7500 160.6000 84.4500 ;
      RECT 0.7000 83.4500 160.6000 83.7500 ;
      RECT 0.0000 82.7500 160.6000 83.4500 ;
      RECT 0.7000 82.4500 160.6000 82.7500 ;
      RECT 0.0000 81.7500 160.6000 82.4500 ;
      RECT 0.7000 81.4500 160.6000 81.7500 ;
      RECT 0.0000 80.7500 160.6000 81.4500 ;
      RECT 0.7000 80.4500 160.6000 80.7500 ;
      RECT 0.0000 79.7500 160.6000 80.4500 ;
      RECT 0.7000 79.4500 160.6000 79.7500 ;
      RECT 0.0000 78.7500 160.6000 79.4500 ;
      RECT 0.7000 78.4500 160.6000 78.7500 ;
      RECT 0.0000 77.7500 160.6000 78.4500 ;
      RECT 0.7000 77.4500 160.6000 77.7500 ;
      RECT 0.0000 76.7500 160.6000 77.4500 ;
      RECT 0.7000 76.4500 160.6000 76.7500 ;
      RECT 0.0000 75.7500 160.6000 76.4500 ;
      RECT 0.7000 75.4500 160.6000 75.7500 ;
      RECT 0.0000 74.7500 160.6000 75.4500 ;
      RECT 0.7000 74.4500 160.6000 74.7500 ;
      RECT 0.0000 73.7500 160.6000 74.4500 ;
      RECT 0.7000 73.4500 160.6000 73.7500 ;
      RECT 0.0000 72.7500 160.6000 73.4500 ;
      RECT 0.7000 72.4500 160.6000 72.7500 ;
      RECT 0.0000 71.7500 160.6000 72.4500 ;
      RECT 0.7000 71.4500 160.6000 71.7500 ;
      RECT 0.0000 70.7500 160.6000 71.4500 ;
      RECT 0.7000 70.4500 160.6000 70.7500 ;
      RECT 0.0000 69.7500 160.6000 70.4500 ;
      RECT 0.7000 69.4500 160.6000 69.7500 ;
      RECT 0.0000 68.7500 160.6000 69.4500 ;
      RECT 0.7000 68.4500 160.6000 68.7500 ;
      RECT 0.0000 67.7500 160.6000 68.4500 ;
      RECT 0.7000 67.4500 160.6000 67.7500 ;
      RECT 0.0000 66.7500 160.6000 67.4500 ;
      RECT 0.7000 66.4500 160.6000 66.7500 ;
      RECT 0.0000 65.7500 160.6000 66.4500 ;
      RECT 0.7000 65.4500 160.6000 65.7500 ;
      RECT 0.0000 64.7500 160.6000 65.4500 ;
      RECT 0.7000 64.4500 160.6000 64.7500 ;
      RECT 0.0000 63.7500 160.6000 64.4500 ;
      RECT 0.7000 63.4500 160.6000 63.7500 ;
      RECT 0.0000 62.7500 160.6000 63.4500 ;
      RECT 0.7000 62.4500 160.6000 62.7500 ;
      RECT 0.0000 61.7500 160.6000 62.4500 ;
      RECT 0.7000 61.4500 160.6000 61.7500 ;
      RECT 0.0000 60.7500 160.6000 61.4500 ;
      RECT 0.7000 60.4500 160.6000 60.7500 ;
      RECT 0.0000 59.7500 160.6000 60.4500 ;
      RECT 0.7000 59.4500 160.6000 59.7500 ;
      RECT 0.0000 58.7500 160.6000 59.4500 ;
      RECT 0.7000 58.4500 160.6000 58.7500 ;
      RECT 0.0000 57.7500 160.6000 58.4500 ;
      RECT 0.7000 57.4500 160.6000 57.7500 ;
      RECT 0.0000 56.7500 160.6000 57.4500 ;
      RECT 0.7000 56.4500 160.6000 56.7500 ;
      RECT 0.0000 55.7500 160.6000 56.4500 ;
      RECT 0.7000 55.4500 160.6000 55.7500 ;
      RECT 0.0000 54.7500 160.6000 55.4500 ;
      RECT 0.7000 54.4500 160.6000 54.7500 ;
      RECT 0.0000 53.7500 160.6000 54.4500 ;
      RECT 0.7000 53.4500 160.6000 53.7500 ;
      RECT 0.0000 52.7500 160.6000 53.4500 ;
      RECT 0.7000 52.4500 160.6000 52.7500 ;
      RECT 0.0000 51.7500 160.6000 52.4500 ;
      RECT 0.7000 51.4500 160.6000 51.7500 ;
      RECT 0.0000 50.7500 160.6000 51.4500 ;
      RECT 0.7000 50.4500 160.6000 50.7500 ;
      RECT 0.0000 49.7500 160.6000 50.4500 ;
      RECT 0.7000 49.4500 160.6000 49.7500 ;
      RECT 0.0000 48.7500 160.6000 49.4500 ;
      RECT 0.7000 48.4500 160.6000 48.7500 ;
      RECT 0.0000 47.7500 160.6000 48.4500 ;
      RECT 0.7000 47.4500 160.6000 47.7500 ;
      RECT 0.0000 46.7500 160.6000 47.4500 ;
      RECT 0.7000 46.4500 160.6000 46.7500 ;
      RECT 0.0000 45.7500 160.6000 46.4500 ;
      RECT 0.7000 45.4500 160.6000 45.7500 ;
      RECT 0.0000 44.7500 160.6000 45.4500 ;
      RECT 0.7000 44.4500 160.6000 44.7500 ;
      RECT 0.0000 43.7500 160.6000 44.4500 ;
      RECT 0.7000 43.4500 160.6000 43.7500 ;
      RECT 0.0000 42.7500 160.6000 43.4500 ;
      RECT 0.7000 42.4500 160.6000 42.7500 ;
      RECT 0.0000 41.7500 160.6000 42.4500 ;
      RECT 0.7000 41.4500 160.6000 41.7500 ;
      RECT 0.0000 40.7500 160.6000 41.4500 ;
      RECT 0.7000 40.4500 160.6000 40.7500 ;
      RECT 0.0000 39.7500 160.6000 40.4500 ;
      RECT 0.7000 39.4500 160.6000 39.7500 ;
      RECT 0.0000 38.7500 160.6000 39.4500 ;
      RECT 0.7000 38.4500 160.6000 38.7500 ;
      RECT 0.0000 37.7500 160.6000 38.4500 ;
      RECT 0.7000 37.4500 160.6000 37.7500 ;
      RECT 0.0000 36.7500 160.6000 37.4500 ;
      RECT 0.7000 36.4500 160.6000 36.7500 ;
      RECT 0.0000 35.7500 160.6000 36.4500 ;
      RECT 0.7000 35.4500 160.6000 35.7500 ;
      RECT 0.0000 34.7500 160.6000 35.4500 ;
      RECT 0.7000 34.4500 160.6000 34.7500 ;
      RECT 0.0000 33.7500 160.6000 34.4500 ;
      RECT 0.7000 33.4500 160.6000 33.7500 ;
      RECT 0.0000 32.7500 160.6000 33.4500 ;
      RECT 0.7000 32.4500 160.6000 32.7500 ;
      RECT 0.0000 31.7500 160.6000 32.4500 ;
      RECT 0.7000 31.4500 160.6000 31.7500 ;
      RECT 0.0000 30.7500 160.6000 31.4500 ;
      RECT 0.7000 30.4500 160.6000 30.7500 ;
      RECT 0.0000 29.7500 160.6000 30.4500 ;
      RECT 0.7000 29.4500 160.6000 29.7500 ;
      RECT 0.0000 28.7500 160.6000 29.4500 ;
      RECT 0.7000 28.4500 160.6000 28.7500 ;
      RECT 0.0000 27.7500 160.6000 28.4500 ;
      RECT 0.7000 27.4500 160.6000 27.7500 ;
      RECT 0.0000 26.7500 160.6000 27.4500 ;
      RECT 0.7000 26.4500 160.6000 26.7500 ;
      RECT 0.0000 25.7500 160.6000 26.4500 ;
      RECT 0.7000 25.4500 160.6000 25.7500 ;
      RECT 0.0000 24.7500 160.6000 25.4500 ;
      RECT 0.7000 24.4500 160.6000 24.7500 ;
      RECT 0.0000 23.7500 160.6000 24.4500 ;
      RECT 0.7000 23.4500 160.6000 23.7500 ;
      RECT 0.0000 22.7500 160.6000 23.4500 ;
      RECT 0.7000 22.4500 160.6000 22.7500 ;
      RECT 0.0000 21.7500 160.6000 22.4500 ;
      RECT 0.7000 21.4500 160.6000 21.7500 ;
      RECT 0.0000 20.7500 160.6000 21.4500 ;
      RECT 0.7000 20.4500 160.6000 20.7500 ;
      RECT 0.0000 19.7500 160.6000 20.4500 ;
      RECT 0.7000 19.4500 160.6000 19.7500 ;
      RECT 0.0000 18.7500 160.6000 19.4500 ;
      RECT 0.7000 18.4500 160.6000 18.7500 ;
      RECT 0.0000 17.7500 160.6000 18.4500 ;
      RECT 0.7000 17.4500 160.6000 17.7500 ;
      RECT 0.0000 16.7500 160.6000 17.4500 ;
      RECT 0.7000 16.4500 160.6000 16.7500 ;
      RECT 0.0000 15.7500 160.6000 16.4500 ;
      RECT 0.7000 15.4500 160.6000 15.7500 ;
      RECT 0.0000 14.7500 160.6000 15.4500 ;
      RECT 0.7000 14.4500 160.6000 14.7500 ;
      RECT 0.0000 0.7600 160.6000 14.4500 ;
      RECT 90.7100 0.0000 160.6000 0.7600 ;
      RECT 89.7100 0.0000 90.2900 0.7600 ;
      RECT 88.7100 0.0000 89.2900 0.7600 ;
      RECT 87.7100 0.0000 88.2900 0.7600 ;
      RECT 86.7100 0.0000 87.2900 0.7600 ;
      RECT 85.7100 0.0000 86.2900 0.7600 ;
      RECT 84.7100 0.0000 85.2900 0.7600 ;
      RECT 83.7100 0.0000 84.2900 0.7600 ;
      RECT 82.7100 0.0000 83.2900 0.7600 ;
      RECT 81.7100 0.0000 82.2900 0.7600 ;
      RECT 80.7100 0.0000 81.2900 0.7600 ;
      RECT 79.7100 0.0000 80.2900 0.7600 ;
      RECT 78.7100 0.0000 79.2900 0.7600 ;
      RECT 77.7100 0.0000 78.2900 0.7600 ;
      RECT 76.7100 0.0000 77.2900 0.7600 ;
      RECT 75.7100 0.0000 76.2900 0.7600 ;
      RECT 74.7100 0.0000 75.2900 0.7600 ;
      RECT 73.7100 0.0000 74.2900 0.7600 ;
      RECT 72.7100 0.0000 73.2900 0.7600 ;
      RECT 71.7100 0.0000 72.2900 0.7600 ;
      RECT 70.7100 0.0000 71.2900 0.7600 ;
      RECT 69.7100 0.0000 70.2900 0.7600 ;
      RECT 0.0000 0.0000 69.2900 0.7600 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 160.6000 158.6000 ;
  END
END mac_8in

END LIBRARY
