/home/linux/ieng6/ee260bwi25/pnataraj/ECE-260B-WI25-Virtuosos/single_core_hierarchical/sram_pnr/sram_w16.lef