##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Mon Mar 17 15:32:17 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO mac_array
  CLASS BLOCK ;
  SIZE 158.6000 BY 155.0000 ;
  FOREIGN mac_array 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 78.9500 158.6000 79.0500 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.0500 154.4800 121.1500 155.0000 ;
    END
  END reset
  PIN in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 154.4800 108.5500 155.0000 ;
    END
  END in[63]
  PIN in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.0500 154.4800 109.1500 155.0000 ;
    END
  END in[62]
  PIN in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.6500 154.4800 109.7500 155.0000 ;
    END
  END in[61]
  PIN in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 108.6500 154.4800 108.7500 155.0000 ;
    END
  END in[60]
  PIN in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.0500 154.4800 100.1500 155.0000 ;
    END
  END in[59]
  PIN in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0500 154.4800 101.1500 155.0000 ;
    END
  END in[58]
  PIN in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.6500 154.4800 100.7500 155.0000 ;
    END
  END in[57]
  PIN in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 109.6500 154.4800 109.7500 155.0000 ;
    END
  END in[56]
  PIN in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 154.4800 74.1500 155.0000 ;
    END
  END in[55]
  PIN in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.0500 154.4800 74.1500 155.0000 ;
    END
  END in[54]
  PIN in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.2500 154.4800 65.3500 155.0000 ;
    END
  END in[53]
  PIN in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 80.1500 0.5200 80.2500 ;
    END
  END in[52]
  PIN in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.6500 154.4800 74.7500 155.0000 ;
    END
  END in[51]
  PIN in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 65.2500 154.4800 65.3500 155.0000 ;
    END
  END in[50]
  PIN in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 78.3500 0.5200 78.4500 ;
    END
  END in[49]
  PIN in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 74.2500 154.4800 74.3500 155.0000 ;
    END
  END in[48]
  PIN in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 154.4800 126.1500 155.0000 ;
    END
  END in[47]
  PIN in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.0500 154.4800 128.1500 155.0000 ;
    END
  END in[46]
  PIN in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.8500 154.4800 135.9500 155.0000 ;
    END
  END in[45]
  PIN in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.6500 154.4800 134.7500 155.0000 ;
    END
  END in[44]
  PIN in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 108.9500 158.6000 109.0500 ;
    END
  END in[43]
  PIN in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 105.3500 158.6000 105.4500 ;
    END
  END in[42]
  PIN in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 134.8500 154.4800 134.9500 155.0000 ;
    END
  END in[41]
  PIN in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 90.9500 158.6000 91.0500 ;
    END
  END in[40]
  PIN in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 29.7500 158.6000 29.8500 ;
    END
  END in[39]
  PIN in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 35.1500 158.6000 35.2500 ;
    END
  END in[38]
  PIN in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 32.3500 158.6000 32.4500 ;
    END
  END in[37]
  PIN in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 39.5500 158.6000 39.6500 ;
    END
  END in[36]
  PIN in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 36.9500 158.6000 37.0500 ;
    END
  END in[35]
  PIN in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 41.5500 158.6000 41.6500 ;
    END
  END in[34]
  PIN in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.6500 0.0000 117.7500 0.5200 ;
    END
  END in[33]
  PIN in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 53.1500 158.6000 53.2500 ;
    END
  END in[32]
  PIN in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 81.1500 158.6000 81.2500 ;
    END
  END in[31]
  PIN in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 91.7500 158.6000 91.8500 ;
    END
  END in[30]
  PIN in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 85.5500 158.6000 85.6500 ;
    END
  END in[29]
  PIN in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.0500 154.4800 83.1500 155.0000 ;
    END
  END in[28]
  PIN in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.0800 90.9500 158.6000 91.0500 ;
    END
  END in[27]
  PIN in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 87.3500 158.6000 87.4500 ;
    END
  END in[26]
  PIN in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 81.9500 158.6000 82.0500 ;
    END
  END in[25]
  PIN in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 80.1500 158.6000 80.2500 ;
    END
  END in[24]
  PIN in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.0500 0.0000 48.1500 0.5200 ;
    END
  END in[23]
  PIN in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 48.0500 0.0000 48.1500 0.5200 ;
    END
  END in[22]
  PIN in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.2500 0.0000 65.3500 0.5200 ;
    END
  END in[21]
  PIN in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 48.0500 0.0000 48.1500 0.5200 ;
    END
  END in[20]
  PIN in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.4500 0.0000 75.5500 0.5200 ;
    END
  END in[19]
  PIN in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.6500 0.0000 74.7500 0.5200 ;
    END
  END in[18]
  PIN in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.0500 0.0000 74.1500 0.5200 ;
    END
  END in[17]
  PIN in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.0500 0.0000 74.1500 0.5200 ;
    END
  END in[16]
  PIN in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.7500 0.5200 56.8500 ;
    END
  END in[15]
  PIN in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.1500 0.5200 53.2500 ;
    END
  END in[14]
  PIN in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.3500 0.5200 69.4500 ;
    END
  END in[13]
  PIN in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 74.7500 0.5200 74.8500 ;
    END
  END in[12]
  PIN in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 62.1500 0.5200 62.2500 ;
    END
  END in[11]
  PIN in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 54.9500 0.5200 55.0500 ;
    END
  END in[10]
  PIN in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 70.3500 0.5200 70.4500 ;
    END
  END in[9]
  PIN in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.9500 0.5200 73.0500 ;
    END
  END in[8]
  PIN in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.4500 0.0000 91.5500 0.5200 ;
    END
  END in[7]
  PIN in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.8500 0.0000 90.9500 0.5200 ;
    END
  END in[6]
  PIN in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.2500 0.0000 109.3500 0.5200 ;
    END
  END in[5]
  PIN in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.0500 0.0000 100.1500 0.5200 ;
    END
  END in[4]
  PIN in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 0.0000 108.5500 0.5200 ;
    END
  END in[3]
  PIN in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.8500 0.0000 112.9500 0.5200 ;
    END
  END in[2]
  PIN in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.2500 0.0000 110.3500 0.5200 ;
    END
  END in[1]
  PIN in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.6500 0.0000 99.7500 0.5200 ;
    END
  END in[0]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 43.7500 158.6000 43.8500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 48.1500 158.6000 48.2500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 76.1500 158.6000 76.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 65.3500 158.6000 65.4500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 66.1500 158.6000 66.2500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 73.3500 158.6000 73.4500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.0800 73.3500 158.6000 73.4500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.6500 154.4800 74.7500 155.0000 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.8500 154.4800 65.9500 155.0000 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.2500 154.4800 57.3500 155.0000 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.8500 154.4800 40.9500 155.0000 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.0500 154.4800 40.1500 155.0000 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 40.0500 154.4800 40.1500 155.0000 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.8500 154.4800 41.9500 155.0000 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 40.0500 154.4800 40.1500 155.0000 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 86.9500 158.6000 87.0500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 83.3500 158.6000 83.4500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 91.3500 158.6000 91.4500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 87.7500 158.6000 87.8500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.0800 87.7500 158.6000 87.8500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 158.0800 80.5500 158.6000 80.6500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M5 ;
        RECT 158.0800 86.9500 158.6000 87.0500 ;
    END
  END out[0]
  PIN fifo_wr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.6500 154.4800 126.7500 155.0000 ;
    END
  END fifo_wr[0]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 125.8500 154.4800 125.9500 155.0000 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M6 ;
        RECT 125.8500 154.4800 125.9500 155.0000 ;
    END
  END inst[0]
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 158.6000 155.0000 ;
    LAYER M2 ;
      RECT 136.0500 154.3800 158.6000 155.0000 ;
      RECT 134.8500 154.3800 135.7500 155.0000 ;
      RECT 128.2500 154.3800 134.5500 155.0000 ;
      RECT 126.8500 154.3800 127.9500 155.0000 ;
      RECT 126.2500 154.3800 126.5500 155.0000 ;
      RECT 121.2500 154.3800 125.9500 155.0000 ;
      RECT 109.8500 154.3800 120.9500 155.0000 ;
      RECT 109.2500 154.3800 109.5500 155.0000 ;
      RECT 108.6500 154.3800 108.9500 155.0000 ;
      RECT 101.2500 154.3800 108.3500 155.0000 ;
      RECT 100.8500 154.3800 100.9500 155.0000 ;
      RECT 100.2500 154.3800 100.5500 155.0000 ;
      RECT 83.2500 154.3800 99.9500 155.0000 ;
      RECT 74.8500 154.3800 82.9500 155.0000 ;
      RECT 74.2500 154.3800 74.5500 155.0000 ;
      RECT 66.0500 154.3800 73.9500 155.0000 ;
      RECT 65.4500 154.3800 65.7500 155.0000 ;
      RECT 57.4500 154.3800 65.1500 155.0000 ;
      RECT 42.0500 154.3800 57.1500 155.0000 ;
      RECT 41.0500 154.3800 41.7500 155.0000 ;
      RECT 40.2500 154.3800 40.7500 155.0000 ;
      RECT 0.0000 154.3800 39.9500 155.0000 ;
      RECT 0.0000 0.6200 158.6000 154.3800 ;
      RECT 117.8500 0.0000 158.6000 0.6200 ;
      RECT 113.0500 0.0000 117.5500 0.6200 ;
      RECT 110.4500 0.0000 112.7500 0.6200 ;
      RECT 109.4500 0.0000 110.1500 0.6200 ;
      RECT 108.6500 0.0000 109.1500 0.6200 ;
      RECT 100.2500 0.0000 108.3500 0.6200 ;
      RECT 99.8500 0.0000 99.9500 0.6200 ;
      RECT 91.6500 0.0000 99.5500 0.6200 ;
      RECT 91.0500 0.0000 91.3500 0.6200 ;
      RECT 75.6500 0.0000 90.7500 0.6200 ;
      RECT 74.8500 0.0000 75.3500 0.6200 ;
      RECT 74.2500 0.0000 74.5500 0.6200 ;
      RECT 65.4500 0.0000 73.9500 0.6200 ;
      RECT 48.2500 0.0000 65.1500 0.6200 ;
      RECT 0.0000 0.0000 47.9500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 109.1500 158.6000 155.0000 ;
      RECT 0.0000 108.8500 157.9800 109.1500 ;
      RECT 0.0000 105.5500 158.6000 108.8500 ;
      RECT 0.0000 105.2500 157.9800 105.5500 ;
      RECT 0.0000 91.9500 158.6000 105.2500 ;
      RECT 0.0000 91.6500 157.9800 91.9500 ;
      RECT 0.0000 91.5500 158.6000 91.6500 ;
      RECT 0.0000 91.2500 157.9800 91.5500 ;
      RECT 0.0000 91.1500 158.6000 91.2500 ;
      RECT 0.0000 90.8500 157.9800 91.1500 ;
      RECT 0.0000 87.9500 158.6000 90.8500 ;
      RECT 0.0000 87.6500 157.9800 87.9500 ;
      RECT 0.0000 87.5500 158.6000 87.6500 ;
      RECT 0.0000 87.2500 157.9800 87.5500 ;
      RECT 0.0000 87.1500 158.6000 87.2500 ;
      RECT 0.0000 86.8500 157.9800 87.1500 ;
      RECT 0.0000 85.7500 158.6000 86.8500 ;
      RECT 0.0000 85.4500 157.9800 85.7500 ;
      RECT 0.0000 83.5500 158.6000 85.4500 ;
      RECT 0.0000 83.2500 157.9800 83.5500 ;
      RECT 0.0000 82.1500 158.6000 83.2500 ;
      RECT 0.0000 81.8500 157.9800 82.1500 ;
      RECT 0.0000 81.3500 158.6000 81.8500 ;
      RECT 0.0000 81.0500 157.9800 81.3500 ;
      RECT 0.0000 80.7500 158.6000 81.0500 ;
      RECT 0.0000 80.4500 157.9800 80.7500 ;
      RECT 0.0000 80.3500 158.6000 80.4500 ;
      RECT 0.6200 80.0500 157.9800 80.3500 ;
      RECT 0.0000 79.1500 158.6000 80.0500 ;
      RECT 0.0000 78.8500 157.9800 79.1500 ;
      RECT 0.0000 78.5500 158.6000 78.8500 ;
      RECT 0.6200 78.2500 158.6000 78.5500 ;
      RECT 0.0000 76.3500 158.6000 78.2500 ;
      RECT 0.0000 76.0500 157.9800 76.3500 ;
      RECT 0.0000 74.9500 158.6000 76.0500 ;
      RECT 0.6200 74.6500 158.6000 74.9500 ;
      RECT 0.0000 73.5500 158.6000 74.6500 ;
      RECT 0.0000 73.2500 157.9800 73.5500 ;
      RECT 0.0000 73.1500 158.6000 73.2500 ;
      RECT 0.6200 72.8500 158.6000 73.1500 ;
      RECT 0.0000 70.5500 158.6000 72.8500 ;
      RECT 0.6200 70.2500 158.6000 70.5500 ;
      RECT 0.0000 69.5500 158.6000 70.2500 ;
      RECT 0.6200 69.2500 158.6000 69.5500 ;
      RECT 0.0000 66.3500 158.6000 69.2500 ;
      RECT 0.0000 66.0500 157.9800 66.3500 ;
      RECT 0.0000 65.5500 158.6000 66.0500 ;
      RECT 0.0000 65.2500 157.9800 65.5500 ;
      RECT 0.0000 62.3500 158.6000 65.2500 ;
      RECT 0.6200 62.0500 158.6000 62.3500 ;
      RECT 0.0000 56.9500 158.6000 62.0500 ;
      RECT 0.6200 56.6500 158.6000 56.9500 ;
      RECT 0.0000 55.1500 158.6000 56.6500 ;
      RECT 0.6200 54.8500 158.6000 55.1500 ;
      RECT 0.0000 53.3500 158.6000 54.8500 ;
      RECT 0.6200 53.0500 157.9800 53.3500 ;
      RECT 0.0000 48.3500 158.6000 53.0500 ;
      RECT 0.0000 48.0500 157.9800 48.3500 ;
      RECT 0.0000 43.9500 158.6000 48.0500 ;
      RECT 0.0000 43.6500 157.9800 43.9500 ;
      RECT 0.0000 41.7500 158.6000 43.6500 ;
      RECT 0.0000 41.4500 157.9800 41.7500 ;
      RECT 0.0000 39.7500 158.6000 41.4500 ;
      RECT 0.0000 39.4500 157.9800 39.7500 ;
      RECT 0.0000 37.1500 158.6000 39.4500 ;
      RECT 0.0000 36.8500 157.9800 37.1500 ;
      RECT 0.0000 35.3500 158.6000 36.8500 ;
      RECT 0.0000 35.0500 157.9800 35.3500 ;
      RECT 0.0000 32.5500 158.6000 35.0500 ;
      RECT 0.0000 32.2500 157.9800 32.5500 ;
      RECT 0.0000 29.9500 158.6000 32.2500 ;
      RECT 0.0000 29.6500 157.9800 29.9500 ;
      RECT 0.0000 0.0000 158.6000 29.6500 ;
    LAYER M4 ;
      RECT 135.0500 154.3800 158.6000 155.0000 ;
      RECT 126.0500 154.3800 134.7500 155.0000 ;
      RECT 109.8500 154.3800 125.7500 155.0000 ;
      RECT 108.8500 154.3800 109.5500 155.0000 ;
      RECT 74.8500 154.3800 108.5500 155.0000 ;
      RECT 74.2500 154.3800 74.5500 155.0000 ;
      RECT 65.4500 154.3800 73.9500 155.0000 ;
      RECT 40.2500 154.3800 65.1500 155.0000 ;
      RECT 0.0000 154.3800 39.9500 155.0000 ;
      RECT 0.0000 0.6200 158.6000 154.3800 ;
      RECT 74.2500 0.0000 158.6000 0.6200 ;
      RECT 48.2500 0.0000 73.9500 0.6200 ;
      RECT 0.0000 0.0000 47.9500 0.6200 ;
    LAYER M5 ;
      RECT 0.0000 91.1500 158.6000 155.0000 ;
      RECT 0.0000 90.8500 157.9800 91.1500 ;
      RECT 0.0000 87.9500 158.6000 90.8500 ;
      RECT 0.0000 87.6500 157.9800 87.9500 ;
      RECT 0.0000 87.1500 158.6000 87.6500 ;
      RECT 0.0000 86.8500 157.9800 87.1500 ;
      RECT 0.0000 73.5500 158.6000 86.8500 ;
      RECT 0.0000 73.2500 157.9800 73.5500 ;
      RECT 0.0000 0.0000 158.6000 73.2500 ;
    LAYER M6 ;
      RECT 126.0500 154.3800 158.6000 155.0000 ;
      RECT 74.4500 154.3800 125.7500 155.0000 ;
      RECT 40.2500 154.3800 74.1500 155.0000 ;
      RECT 0.0000 154.3800 39.9500 155.0000 ;
      RECT 0.0000 0.6200 158.6000 154.3800 ;
      RECT 48.2500 0.0000 158.6000 0.6200 ;
      RECT 0.0000 0.0000 47.9500 0.6200 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 158.6000 155.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 158.6000 155.0000 ;
  END
END mac_array

END LIBRARY
