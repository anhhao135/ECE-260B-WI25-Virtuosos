##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 15 15:47:46 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 286.4000 BY 284.8000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.9500 0.6000 20.0500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.4500 0.0000 92.5500 0.6000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.2500 0.0000 93.3500 0.6000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 0.0000 94.1500 0.6000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 0.0000 94.9500 0.6000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.6500 0.0000 95.7500 0.6000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.4500 0.0000 96.5500 0.6000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.2500 0.0000 97.3500 0.6000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 0.0000 98.1500 0.6000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 0.0000 98.9500 0.6000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.6500 0.0000 99.7500 0.6000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.4500 0.0000 100.5500 0.6000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.2500 0.0000 101.3500 0.6000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 0.0000 102.1500 0.6000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 0.0000 102.9500 0.6000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.6500 0.0000 103.7500 0.6000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4500 0.0000 104.5500 0.6000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.2500 0.0000 105.3500 0.6000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 0.0000 106.1500 0.6000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 0.0000 106.9500 0.6000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.6500 0.0000 107.7500 0.6000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 0.0000 108.5500 0.6000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.2500 0.0000 109.3500 0.6000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 0.0000 110.1500 0.6000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 0.0000 110.9500 0.6000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.6500 0.0000 111.7500 0.6000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.4500 0.0000 112.5500 0.6000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.2500 0.0000 113.3500 0.6000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.0500 0.0000 114.1500 0.6000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 0.0000 114.9500 0.6000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.6500 0.0000 115.7500 0.6000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.4500 0.0000 116.5500 0.6000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.2500 0.0000 117.3500 0.6000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.0500 0.0000 118.1500 0.6000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 0.0000 118.9500 0.6000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.6500 0.0000 119.7500 0.6000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.4500 0.0000 120.5500 0.6000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.2500 0.0000 121.3500 0.6000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.0500 0.0000 122.1500 0.6000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 0.0000 122.9500 0.6000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.6500 0.0000 123.7500 0.6000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.4500 0.0000 124.5500 0.6000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.2500 0.0000 125.3500 0.6000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 0.0000 126.1500 0.6000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 0.0000 126.9500 0.6000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.6500 0.0000 127.7500 0.6000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.4500 0.0000 128.5500 0.6000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.2500 0.0000 129.3500 0.6000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.0500 0.0000 130.1500 0.6000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 0.0000 130.9500 0.6000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.6500 0.0000 131.7500 0.6000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.4500 0.0000 132.5500 0.6000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.2500 0.0000 133.3500 0.6000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 0.0000 134.1500 0.6000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 0.0000 134.9500 0.6000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.6500 0.0000 135.7500 0.6000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.4500 0.0000 136.5500 0.6000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.2500 0.0000 137.3500 0.6000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.0500 0.0000 138.1500 0.6000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 0.0000 138.9500 0.6000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.6500 0.0000 139.7500 0.6000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.4500 0.0000 140.5500 0.6000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.2500 0.0000 141.3500 0.6000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.0500 0.0000 142.1500 0.6000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 0.0000 142.9500 0.6000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.6500 0.0000 143.7500 0.6000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.4500 0.0000 144.5500 0.6000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.2500 0.0000 145.3500 0.6000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.0500 0.0000 146.1500 0.6000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 0.0000 146.9500 0.6000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.6500 0.0000 147.7500 0.6000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.4500 0.0000 148.5500 0.6000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.2500 0.0000 149.3500 0.6000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.0500 0.0000 150.1500 0.6000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 0.0000 150.9500 0.6000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.6500 0.0000 151.7500 0.6000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.4500 0.0000 152.5500 0.6000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.2500 0.0000 153.3500 0.6000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.0500 0.0000 154.1500 0.6000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 0.0000 154.9500 0.6000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.6500 0.0000 155.7500 0.6000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.4500 0.0000 156.5500 0.6000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.2500 0.0000 157.3500 0.6000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.0500 0.0000 158.1500 0.6000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 0.0000 158.9500 0.6000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.6500 0.0000 159.7500 0.6000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.4500 0.0000 160.5500 0.6000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.2500 0.0000 161.3500 0.6000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.0500 0.0000 162.1500 0.6000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 0.0000 162.9500 0.6000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.6500 0.0000 163.7500 0.6000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.4500 0.0000 164.5500 0.6000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.2500 0.0000 165.3500 0.6000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.0500 0.0000 166.1500 0.6000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 0.0000 166.9500 0.6000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.6500 0.0000 167.7500 0.6000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.4500 0.0000 168.5500 0.6000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.2500 0.0000 169.3500 0.6000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.0500 0.0000 170.1500 0.6000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.8500 0.0000 170.9500 0.6000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.6500 0.0000 171.7500 0.6000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.4500 0.0000 172.5500 0.6000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.2500 0.0000 173.3500 0.6000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.0500 0.0000 174.1500 0.6000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.8500 0.0000 174.9500 0.6000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.6500 0.0000 175.7500 0.6000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.4500 0.0000 176.5500 0.6000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.2500 0.0000 177.3500 0.6000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.0500 0.0000 178.1500 0.6000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.8500 0.0000 178.9500 0.6000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.6500 0.0000 179.7500 0.6000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.4500 0.0000 180.5500 0.6000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.2500 0.0000 181.3500 0.6000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.0500 0.0000 182.1500 0.6000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.8500 0.0000 182.9500 0.6000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.6500 0.0000 183.7500 0.6000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.4500 0.0000 184.5500 0.6000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.2500 0.0000 185.3500 0.6000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.0500 0.0000 186.1500 0.6000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.8500 0.0000 186.9500 0.6000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.6500 0.0000 187.7500 0.6000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.4500 0.0000 188.5500 0.6000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.2500 0.0000 189.3500 0.6000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.0500 0.0000 190.1500 0.6000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.8500 0.0000 190.9500 0.6000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.6500 0.0000 191.7500 0.6000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.4500 0.0000 192.5500 0.6000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.2500 0.0000 193.3500 0.6000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.0500 0.0000 194.1500 0.6000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.4500 284.2000 92.5500 284.8000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.2500 284.2000 93.3500 284.8000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.0500 284.2000 94.1500 284.8000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.8500 284.2000 94.9500 284.8000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.6500 284.2000 95.7500 284.8000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.4500 284.2000 96.5500 284.8000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.2500 284.2000 97.3500 284.8000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.0500 284.2000 98.1500 284.8000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.8500 284.2000 98.9500 284.8000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.6500 284.2000 99.7500 284.8000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.4500 284.2000 100.5500 284.8000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.2500 284.2000 101.3500 284.8000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.0500 284.2000 102.1500 284.8000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.8500 284.2000 102.9500 284.8000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.6500 284.2000 103.7500 284.8000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.4500 284.2000 104.5500 284.8000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.2500 284.2000 105.3500 284.8000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.0500 284.2000 106.1500 284.8000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.8500 284.2000 106.9500 284.8000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.6500 284.2000 107.7500 284.8000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.4500 284.2000 108.5500 284.8000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.2500 284.2000 109.3500 284.8000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.0500 284.2000 110.1500 284.8000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.8500 284.2000 110.9500 284.8000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.6500 284.2000 111.7500 284.8000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.4500 284.2000 112.5500 284.8000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.2500 284.2000 113.3500 284.8000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.0500 284.2000 114.1500 284.8000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.8500 284.2000 114.9500 284.8000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.6500 284.2000 115.7500 284.8000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.4500 284.2000 116.5500 284.8000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.2500 284.2000 117.3500 284.8000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.0500 284.2000 118.1500 284.8000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.8500 284.2000 118.9500 284.8000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.6500 284.2000 119.7500 284.8000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.4500 284.2000 120.5500 284.8000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.2500 284.2000 121.3500 284.8000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.0500 284.2000 122.1500 284.8000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.8500 284.2000 122.9500 284.8000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.6500 284.2000 123.7500 284.8000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.4500 284.2000 124.5500 284.8000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.2500 284.2000 125.3500 284.8000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.0500 284.2000 126.1500 284.8000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.8500 284.2000 126.9500 284.8000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.6500 284.2000 127.7500 284.8000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.4500 284.2000 128.5500 284.8000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.2500 284.2000 129.3500 284.8000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.0500 284.2000 130.1500 284.8000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.8500 284.2000 130.9500 284.8000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.6500 284.2000 131.7500 284.8000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.4500 284.2000 132.5500 284.8000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.2500 284.2000 133.3500 284.8000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 284.2000 134.1500 284.8000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.8500 284.2000 134.9500 284.8000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.6500 284.2000 135.7500 284.8000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.4500 284.2000 136.5500 284.8000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.2500 284.2000 137.3500 284.8000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.0500 284.2000 138.1500 284.8000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.8500 284.2000 138.9500 284.8000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.6500 284.2000 139.7500 284.8000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.4500 284.2000 140.5500 284.8000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.2500 284.2000 141.3500 284.8000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.0500 284.2000 142.1500 284.8000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.8500 284.2000 142.9500 284.8000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.6500 284.2000 143.7500 284.8000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.4500 284.2000 144.5500 284.8000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.2500 284.2000 145.3500 284.8000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.0500 284.2000 146.1500 284.8000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.8500 284.2000 146.9500 284.8000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.6500 284.2000 147.7500 284.8000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.4500 284.2000 148.5500 284.8000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.2500 284.2000 149.3500 284.8000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.0500 284.2000 150.1500 284.8000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.8500 284.2000 150.9500 284.8000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.6500 284.2000 151.7500 284.8000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.4500 284.2000 152.5500 284.8000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.2500 284.2000 153.3500 284.8000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.0500 284.2000 154.1500 284.8000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.8500 284.2000 154.9500 284.8000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.6500 284.2000 155.7500 284.8000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.4500 284.2000 156.5500 284.8000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.2500 284.2000 157.3500 284.8000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.0500 284.2000 158.1500 284.8000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.8500 284.2000 158.9500 284.8000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.6500 284.2000 159.7500 284.8000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.4500 284.2000 160.5500 284.8000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.2500 284.2000 161.3500 284.8000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.0500 284.2000 162.1500 284.8000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.8500 284.2000 162.9500 284.8000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.6500 284.2000 163.7500 284.8000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.4500 284.2000 164.5500 284.8000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.2500 284.2000 165.3500 284.8000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.0500 284.2000 166.1500 284.8000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.8500 284.2000 166.9500 284.8000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.6500 284.2000 167.7500 284.8000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.4500 284.2000 168.5500 284.8000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.2500 284.2000 169.3500 284.8000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.0500 284.2000 170.1500 284.8000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.8500 284.2000 170.9500 284.8000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.6500 284.2000 171.7500 284.8000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.4500 284.2000 172.5500 284.8000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.2500 284.2000 173.3500 284.8000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.0500 284.2000 174.1500 284.8000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 174.8500 284.2000 174.9500 284.8000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.6500 284.2000 175.7500 284.8000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.4500 284.2000 176.5500 284.8000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.2500 284.2000 177.3500 284.8000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.0500 284.2000 178.1500 284.8000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.8500 284.2000 178.9500 284.8000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.6500 284.2000 179.7500 284.8000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.4500 284.2000 180.5500 284.8000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.2500 284.2000 181.3500 284.8000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.0500 284.2000 182.1500 284.8000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.8500 284.2000 182.9500 284.8000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.6500 284.2000 183.7500 284.8000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.4500 284.2000 184.5500 284.8000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.2500 284.2000 185.3500 284.8000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.0500 284.2000 186.1500 284.8000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.8500 284.2000 186.9500 284.8000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.6500 284.2000 187.7500 284.8000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.4500 284.2000 188.5500 284.8000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.2500 284.2000 189.3500 284.8000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.0500 284.2000 190.1500 284.8000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.8500 284.2000 190.9500 284.8000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.6500 284.2000 191.7500 284.8000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.4500 284.2000 192.5500 284.8000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.2500 284.2000 193.3500 284.8000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.0500 284.2000 194.1500 284.8000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 19.1500 0.6000 19.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 20.7500 0.6000 20.8500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 18.3500 0.6000 18.4500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.5500 0.6000 17.6500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 16.7500 0.6000 16.8500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 15.9500 0.6000 16.0500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 28.0000 20.0000 30.0000 264.8000 ;
        RECT 54.2650 20.0000 56.2650 264.8000 ;
        RECT 80.5300 20.0000 82.5300 264.8000 ;
        RECT 106.7950 20.0000 108.7950 264.8000 ;
        RECT 133.0600 20.0000 135.0600 264.8000 ;
        RECT 159.3250 20.0000 161.3250 264.8000 ;
        RECT 185.5900 20.0000 187.5900 264.8000 ;
        RECT 211.8550 20.0000 213.8550 264.8000 ;
        RECT 238.1200 20.0000 240.1200 264.8000 ;
        RECT 264.3850 20.0000 266.3850 264.8000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 20.0000 20.0000 22.0000 264.8000 ;
        RECT 46.2650 20.0000 48.2650 264.8000 ;
        RECT 72.5300 20.0000 74.5300 264.8000 ;
        RECT 98.7950 20.0000 100.7950 264.8000 ;
        RECT 125.0600 20.0000 127.0600 264.8000 ;
        RECT 151.3250 20.0000 153.3250 264.8000 ;
        RECT 177.5900 20.0000 179.5900 264.8000 ;
        RECT 203.8550 20.0000 205.8550 264.8000 ;
        RECT 230.1200 20.0000 232.1200 264.8000 ;
        RECT 256.3850 20.0000 258.3850 264.8000 ;
        RECT 20.0000 19.8350 22.0000 20.1650 ;
        RECT 46.2650 19.8350 48.2650 20.1650 ;
        RECT 72.5300 19.8350 74.5300 20.1650 ;
        RECT 98.7950 19.8350 100.7950 20.1650 ;
        RECT 125.0600 19.8350 127.0600 20.1650 ;
        RECT 177.5900 19.8350 179.5900 20.1650 ;
        RECT 151.3250 19.8350 153.3250 20.1650 ;
        RECT 203.8550 19.8350 205.8550 20.1650 ;
        RECT 230.1200 19.8350 232.1200 20.1650 ;
        RECT 256.3850 19.8350 258.3850 20.1650 ;
        RECT 20.0000 264.6350 22.0000 264.9650 ;
        RECT 46.2650 264.6350 48.2650 264.9650 ;
        RECT 72.5300 264.6350 74.5300 264.9650 ;
        RECT 98.7950 264.6350 100.7950 264.9650 ;
        RECT 125.0600 264.6350 127.0600 264.9650 ;
        RECT 177.5900 264.6350 179.5900 264.9650 ;
        RECT 151.3250 264.6350 153.3250 264.9650 ;
        RECT 203.8550 264.6350 205.8550 264.9650 ;
        RECT 230.1200 264.6350 232.1200 264.9650 ;
        RECT 256.3850 264.6350 258.3850 264.9650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 286.4000 284.8000 ;
    LAYER M2 ;
      RECT 194.2500 284.1000 286.4000 284.8000 ;
      RECT 193.4500 284.1000 193.9500 284.8000 ;
      RECT 192.6500 284.1000 193.1500 284.8000 ;
      RECT 191.8500 284.1000 192.3500 284.8000 ;
      RECT 191.0500 284.1000 191.5500 284.8000 ;
      RECT 190.2500 284.1000 190.7500 284.8000 ;
      RECT 189.4500 284.1000 189.9500 284.8000 ;
      RECT 188.6500 284.1000 189.1500 284.8000 ;
      RECT 187.8500 284.1000 188.3500 284.8000 ;
      RECT 187.0500 284.1000 187.5500 284.8000 ;
      RECT 186.2500 284.1000 186.7500 284.8000 ;
      RECT 185.4500 284.1000 185.9500 284.8000 ;
      RECT 184.6500 284.1000 185.1500 284.8000 ;
      RECT 183.8500 284.1000 184.3500 284.8000 ;
      RECT 183.0500 284.1000 183.5500 284.8000 ;
      RECT 182.2500 284.1000 182.7500 284.8000 ;
      RECT 181.4500 284.1000 181.9500 284.8000 ;
      RECT 180.6500 284.1000 181.1500 284.8000 ;
      RECT 179.8500 284.1000 180.3500 284.8000 ;
      RECT 179.0500 284.1000 179.5500 284.8000 ;
      RECT 178.2500 284.1000 178.7500 284.8000 ;
      RECT 177.4500 284.1000 177.9500 284.8000 ;
      RECT 176.6500 284.1000 177.1500 284.8000 ;
      RECT 175.8500 284.1000 176.3500 284.8000 ;
      RECT 175.0500 284.1000 175.5500 284.8000 ;
      RECT 174.2500 284.1000 174.7500 284.8000 ;
      RECT 173.4500 284.1000 173.9500 284.8000 ;
      RECT 172.6500 284.1000 173.1500 284.8000 ;
      RECT 171.8500 284.1000 172.3500 284.8000 ;
      RECT 171.0500 284.1000 171.5500 284.8000 ;
      RECT 170.2500 284.1000 170.7500 284.8000 ;
      RECT 169.4500 284.1000 169.9500 284.8000 ;
      RECT 168.6500 284.1000 169.1500 284.8000 ;
      RECT 167.8500 284.1000 168.3500 284.8000 ;
      RECT 167.0500 284.1000 167.5500 284.8000 ;
      RECT 166.2500 284.1000 166.7500 284.8000 ;
      RECT 165.4500 284.1000 165.9500 284.8000 ;
      RECT 164.6500 284.1000 165.1500 284.8000 ;
      RECT 163.8500 284.1000 164.3500 284.8000 ;
      RECT 163.0500 284.1000 163.5500 284.8000 ;
      RECT 162.2500 284.1000 162.7500 284.8000 ;
      RECT 161.4500 284.1000 161.9500 284.8000 ;
      RECT 160.6500 284.1000 161.1500 284.8000 ;
      RECT 159.8500 284.1000 160.3500 284.8000 ;
      RECT 159.0500 284.1000 159.5500 284.8000 ;
      RECT 158.2500 284.1000 158.7500 284.8000 ;
      RECT 157.4500 284.1000 157.9500 284.8000 ;
      RECT 156.6500 284.1000 157.1500 284.8000 ;
      RECT 155.8500 284.1000 156.3500 284.8000 ;
      RECT 155.0500 284.1000 155.5500 284.8000 ;
      RECT 154.2500 284.1000 154.7500 284.8000 ;
      RECT 153.4500 284.1000 153.9500 284.8000 ;
      RECT 152.6500 284.1000 153.1500 284.8000 ;
      RECT 151.8500 284.1000 152.3500 284.8000 ;
      RECT 151.0500 284.1000 151.5500 284.8000 ;
      RECT 150.2500 284.1000 150.7500 284.8000 ;
      RECT 149.4500 284.1000 149.9500 284.8000 ;
      RECT 148.6500 284.1000 149.1500 284.8000 ;
      RECT 147.8500 284.1000 148.3500 284.8000 ;
      RECT 147.0500 284.1000 147.5500 284.8000 ;
      RECT 146.2500 284.1000 146.7500 284.8000 ;
      RECT 145.4500 284.1000 145.9500 284.8000 ;
      RECT 144.6500 284.1000 145.1500 284.8000 ;
      RECT 143.8500 284.1000 144.3500 284.8000 ;
      RECT 143.0500 284.1000 143.5500 284.8000 ;
      RECT 142.2500 284.1000 142.7500 284.8000 ;
      RECT 141.4500 284.1000 141.9500 284.8000 ;
      RECT 140.6500 284.1000 141.1500 284.8000 ;
      RECT 139.8500 284.1000 140.3500 284.8000 ;
      RECT 139.0500 284.1000 139.5500 284.8000 ;
      RECT 138.2500 284.1000 138.7500 284.8000 ;
      RECT 137.4500 284.1000 137.9500 284.8000 ;
      RECT 136.6500 284.1000 137.1500 284.8000 ;
      RECT 135.8500 284.1000 136.3500 284.8000 ;
      RECT 135.0500 284.1000 135.5500 284.8000 ;
      RECT 134.2500 284.1000 134.7500 284.8000 ;
      RECT 133.4500 284.1000 133.9500 284.8000 ;
      RECT 132.6500 284.1000 133.1500 284.8000 ;
      RECT 131.8500 284.1000 132.3500 284.8000 ;
      RECT 131.0500 284.1000 131.5500 284.8000 ;
      RECT 130.2500 284.1000 130.7500 284.8000 ;
      RECT 129.4500 284.1000 129.9500 284.8000 ;
      RECT 128.6500 284.1000 129.1500 284.8000 ;
      RECT 127.8500 284.1000 128.3500 284.8000 ;
      RECT 127.0500 284.1000 127.5500 284.8000 ;
      RECT 126.2500 284.1000 126.7500 284.8000 ;
      RECT 125.4500 284.1000 125.9500 284.8000 ;
      RECT 124.6500 284.1000 125.1500 284.8000 ;
      RECT 123.8500 284.1000 124.3500 284.8000 ;
      RECT 123.0500 284.1000 123.5500 284.8000 ;
      RECT 122.2500 284.1000 122.7500 284.8000 ;
      RECT 121.4500 284.1000 121.9500 284.8000 ;
      RECT 120.6500 284.1000 121.1500 284.8000 ;
      RECT 119.8500 284.1000 120.3500 284.8000 ;
      RECT 119.0500 284.1000 119.5500 284.8000 ;
      RECT 118.2500 284.1000 118.7500 284.8000 ;
      RECT 117.4500 284.1000 117.9500 284.8000 ;
      RECT 116.6500 284.1000 117.1500 284.8000 ;
      RECT 115.8500 284.1000 116.3500 284.8000 ;
      RECT 115.0500 284.1000 115.5500 284.8000 ;
      RECT 114.2500 284.1000 114.7500 284.8000 ;
      RECT 113.4500 284.1000 113.9500 284.8000 ;
      RECT 112.6500 284.1000 113.1500 284.8000 ;
      RECT 111.8500 284.1000 112.3500 284.8000 ;
      RECT 111.0500 284.1000 111.5500 284.8000 ;
      RECT 110.2500 284.1000 110.7500 284.8000 ;
      RECT 109.4500 284.1000 109.9500 284.8000 ;
      RECT 108.6500 284.1000 109.1500 284.8000 ;
      RECT 107.8500 284.1000 108.3500 284.8000 ;
      RECT 107.0500 284.1000 107.5500 284.8000 ;
      RECT 106.2500 284.1000 106.7500 284.8000 ;
      RECT 105.4500 284.1000 105.9500 284.8000 ;
      RECT 104.6500 284.1000 105.1500 284.8000 ;
      RECT 103.8500 284.1000 104.3500 284.8000 ;
      RECT 103.0500 284.1000 103.5500 284.8000 ;
      RECT 102.2500 284.1000 102.7500 284.8000 ;
      RECT 101.4500 284.1000 101.9500 284.8000 ;
      RECT 100.6500 284.1000 101.1500 284.8000 ;
      RECT 99.8500 284.1000 100.3500 284.8000 ;
      RECT 99.0500 284.1000 99.5500 284.8000 ;
      RECT 98.2500 284.1000 98.7500 284.8000 ;
      RECT 97.4500 284.1000 97.9500 284.8000 ;
      RECT 96.6500 284.1000 97.1500 284.8000 ;
      RECT 95.8500 284.1000 96.3500 284.8000 ;
      RECT 95.0500 284.1000 95.5500 284.8000 ;
      RECT 94.2500 284.1000 94.7500 284.8000 ;
      RECT 93.4500 284.1000 93.9500 284.8000 ;
      RECT 92.6500 284.1000 93.1500 284.8000 ;
      RECT 0.0000 284.1000 92.3500 284.8000 ;
      RECT 0.0000 0.7000 286.4000 284.1000 ;
      RECT 194.2500 0.0000 286.4000 0.7000 ;
      RECT 193.4500 0.0000 193.9500 0.7000 ;
      RECT 192.6500 0.0000 193.1500 0.7000 ;
      RECT 191.8500 0.0000 192.3500 0.7000 ;
      RECT 191.0500 0.0000 191.5500 0.7000 ;
      RECT 190.2500 0.0000 190.7500 0.7000 ;
      RECT 189.4500 0.0000 189.9500 0.7000 ;
      RECT 188.6500 0.0000 189.1500 0.7000 ;
      RECT 187.8500 0.0000 188.3500 0.7000 ;
      RECT 187.0500 0.0000 187.5500 0.7000 ;
      RECT 186.2500 0.0000 186.7500 0.7000 ;
      RECT 185.4500 0.0000 185.9500 0.7000 ;
      RECT 184.6500 0.0000 185.1500 0.7000 ;
      RECT 183.8500 0.0000 184.3500 0.7000 ;
      RECT 183.0500 0.0000 183.5500 0.7000 ;
      RECT 182.2500 0.0000 182.7500 0.7000 ;
      RECT 181.4500 0.0000 181.9500 0.7000 ;
      RECT 180.6500 0.0000 181.1500 0.7000 ;
      RECT 179.8500 0.0000 180.3500 0.7000 ;
      RECT 179.0500 0.0000 179.5500 0.7000 ;
      RECT 178.2500 0.0000 178.7500 0.7000 ;
      RECT 177.4500 0.0000 177.9500 0.7000 ;
      RECT 176.6500 0.0000 177.1500 0.7000 ;
      RECT 175.8500 0.0000 176.3500 0.7000 ;
      RECT 175.0500 0.0000 175.5500 0.7000 ;
      RECT 174.2500 0.0000 174.7500 0.7000 ;
      RECT 173.4500 0.0000 173.9500 0.7000 ;
      RECT 172.6500 0.0000 173.1500 0.7000 ;
      RECT 171.8500 0.0000 172.3500 0.7000 ;
      RECT 171.0500 0.0000 171.5500 0.7000 ;
      RECT 170.2500 0.0000 170.7500 0.7000 ;
      RECT 169.4500 0.0000 169.9500 0.7000 ;
      RECT 168.6500 0.0000 169.1500 0.7000 ;
      RECT 167.8500 0.0000 168.3500 0.7000 ;
      RECT 167.0500 0.0000 167.5500 0.7000 ;
      RECT 166.2500 0.0000 166.7500 0.7000 ;
      RECT 165.4500 0.0000 165.9500 0.7000 ;
      RECT 164.6500 0.0000 165.1500 0.7000 ;
      RECT 163.8500 0.0000 164.3500 0.7000 ;
      RECT 163.0500 0.0000 163.5500 0.7000 ;
      RECT 162.2500 0.0000 162.7500 0.7000 ;
      RECT 161.4500 0.0000 161.9500 0.7000 ;
      RECT 160.6500 0.0000 161.1500 0.7000 ;
      RECT 159.8500 0.0000 160.3500 0.7000 ;
      RECT 159.0500 0.0000 159.5500 0.7000 ;
      RECT 158.2500 0.0000 158.7500 0.7000 ;
      RECT 157.4500 0.0000 157.9500 0.7000 ;
      RECT 156.6500 0.0000 157.1500 0.7000 ;
      RECT 155.8500 0.0000 156.3500 0.7000 ;
      RECT 155.0500 0.0000 155.5500 0.7000 ;
      RECT 154.2500 0.0000 154.7500 0.7000 ;
      RECT 153.4500 0.0000 153.9500 0.7000 ;
      RECT 152.6500 0.0000 153.1500 0.7000 ;
      RECT 151.8500 0.0000 152.3500 0.7000 ;
      RECT 151.0500 0.0000 151.5500 0.7000 ;
      RECT 150.2500 0.0000 150.7500 0.7000 ;
      RECT 149.4500 0.0000 149.9500 0.7000 ;
      RECT 148.6500 0.0000 149.1500 0.7000 ;
      RECT 147.8500 0.0000 148.3500 0.7000 ;
      RECT 147.0500 0.0000 147.5500 0.7000 ;
      RECT 146.2500 0.0000 146.7500 0.7000 ;
      RECT 145.4500 0.0000 145.9500 0.7000 ;
      RECT 144.6500 0.0000 145.1500 0.7000 ;
      RECT 143.8500 0.0000 144.3500 0.7000 ;
      RECT 143.0500 0.0000 143.5500 0.7000 ;
      RECT 142.2500 0.0000 142.7500 0.7000 ;
      RECT 141.4500 0.0000 141.9500 0.7000 ;
      RECT 140.6500 0.0000 141.1500 0.7000 ;
      RECT 139.8500 0.0000 140.3500 0.7000 ;
      RECT 139.0500 0.0000 139.5500 0.7000 ;
      RECT 138.2500 0.0000 138.7500 0.7000 ;
      RECT 137.4500 0.0000 137.9500 0.7000 ;
      RECT 136.6500 0.0000 137.1500 0.7000 ;
      RECT 135.8500 0.0000 136.3500 0.7000 ;
      RECT 135.0500 0.0000 135.5500 0.7000 ;
      RECT 134.2500 0.0000 134.7500 0.7000 ;
      RECT 133.4500 0.0000 133.9500 0.7000 ;
      RECT 132.6500 0.0000 133.1500 0.7000 ;
      RECT 131.8500 0.0000 132.3500 0.7000 ;
      RECT 131.0500 0.0000 131.5500 0.7000 ;
      RECT 130.2500 0.0000 130.7500 0.7000 ;
      RECT 129.4500 0.0000 129.9500 0.7000 ;
      RECT 128.6500 0.0000 129.1500 0.7000 ;
      RECT 127.8500 0.0000 128.3500 0.7000 ;
      RECT 127.0500 0.0000 127.5500 0.7000 ;
      RECT 126.2500 0.0000 126.7500 0.7000 ;
      RECT 125.4500 0.0000 125.9500 0.7000 ;
      RECT 124.6500 0.0000 125.1500 0.7000 ;
      RECT 123.8500 0.0000 124.3500 0.7000 ;
      RECT 123.0500 0.0000 123.5500 0.7000 ;
      RECT 122.2500 0.0000 122.7500 0.7000 ;
      RECT 121.4500 0.0000 121.9500 0.7000 ;
      RECT 120.6500 0.0000 121.1500 0.7000 ;
      RECT 119.8500 0.0000 120.3500 0.7000 ;
      RECT 119.0500 0.0000 119.5500 0.7000 ;
      RECT 118.2500 0.0000 118.7500 0.7000 ;
      RECT 117.4500 0.0000 117.9500 0.7000 ;
      RECT 116.6500 0.0000 117.1500 0.7000 ;
      RECT 115.8500 0.0000 116.3500 0.7000 ;
      RECT 115.0500 0.0000 115.5500 0.7000 ;
      RECT 114.2500 0.0000 114.7500 0.7000 ;
      RECT 113.4500 0.0000 113.9500 0.7000 ;
      RECT 112.6500 0.0000 113.1500 0.7000 ;
      RECT 111.8500 0.0000 112.3500 0.7000 ;
      RECT 111.0500 0.0000 111.5500 0.7000 ;
      RECT 110.2500 0.0000 110.7500 0.7000 ;
      RECT 109.4500 0.0000 109.9500 0.7000 ;
      RECT 108.6500 0.0000 109.1500 0.7000 ;
      RECT 107.8500 0.0000 108.3500 0.7000 ;
      RECT 107.0500 0.0000 107.5500 0.7000 ;
      RECT 106.2500 0.0000 106.7500 0.7000 ;
      RECT 105.4500 0.0000 105.9500 0.7000 ;
      RECT 104.6500 0.0000 105.1500 0.7000 ;
      RECT 103.8500 0.0000 104.3500 0.7000 ;
      RECT 103.0500 0.0000 103.5500 0.7000 ;
      RECT 102.2500 0.0000 102.7500 0.7000 ;
      RECT 101.4500 0.0000 101.9500 0.7000 ;
      RECT 100.6500 0.0000 101.1500 0.7000 ;
      RECT 99.8500 0.0000 100.3500 0.7000 ;
      RECT 99.0500 0.0000 99.5500 0.7000 ;
      RECT 98.2500 0.0000 98.7500 0.7000 ;
      RECT 97.4500 0.0000 97.9500 0.7000 ;
      RECT 96.6500 0.0000 97.1500 0.7000 ;
      RECT 95.8500 0.0000 96.3500 0.7000 ;
      RECT 95.0500 0.0000 95.5500 0.7000 ;
      RECT 94.2500 0.0000 94.7500 0.7000 ;
      RECT 93.4500 0.0000 93.9500 0.7000 ;
      RECT 92.6500 0.0000 93.1500 0.7000 ;
      RECT 0.0000 0.0000 92.3500 0.7000 ;
    LAYER M3 ;
      RECT 0.0000 20.9500 286.4000 284.8000 ;
      RECT 0.7000 20.6500 286.4000 20.9500 ;
      RECT 0.0000 20.1500 286.4000 20.6500 ;
      RECT 0.7000 19.8500 286.4000 20.1500 ;
      RECT 0.0000 19.3500 286.4000 19.8500 ;
      RECT 0.7000 19.0500 286.4000 19.3500 ;
      RECT 0.0000 18.5500 286.4000 19.0500 ;
      RECT 0.7000 18.2500 286.4000 18.5500 ;
      RECT 0.0000 17.7500 286.4000 18.2500 ;
      RECT 0.7000 17.4500 286.4000 17.7500 ;
      RECT 0.0000 16.9500 286.4000 17.4500 ;
      RECT 0.7000 16.6500 286.4000 16.9500 ;
      RECT 0.0000 16.1500 286.4000 16.6500 ;
      RECT 0.7000 15.8500 286.4000 16.1500 ;
      RECT 0.0000 0.0000 286.4000 15.8500 ;
    LAYER M4 ;
      RECT 0.0000 265.4650 286.4000 284.8000 ;
      RECT 258.8850 265.3000 286.4000 265.4650 ;
      RECT 232.6200 265.3000 255.8850 265.4650 ;
      RECT 206.3550 265.3000 229.6200 265.4650 ;
      RECT 180.0900 265.3000 203.3550 265.4650 ;
      RECT 153.8250 265.3000 177.0900 265.4650 ;
      RECT 127.5600 265.3000 150.8250 265.4650 ;
      RECT 101.2950 265.3000 124.5600 265.4650 ;
      RECT 75.0300 265.3000 98.2950 265.4650 ;
      RECT 48.7650 265.3000 72.0300 265.4650 ;
      RECT 22.5000 265.3000 45.7650 265.4650 ;
      RECT 266.8850 19.5000 286.4000 265.3000 ;
      RECT 258.8850 19.5000 263.8850 265.3000 ;
      RECT 240.6200 19.5000 255.8850 265.3000 ;
      RECT 232.6200 19.5000 237.6200 265.3000 ;
      RECT 214.3550 19.5000 229.6200 265.3000 ;
      RECT 206.3550 19.5000 211.3550 265.3000 ;
      RECT 188.0900 19.5000 203.3550 265.3000 ;
      RECT 180.0900 19.5000 185.0900 265.3000 ;
      RECT 161.8250 19.5000 177.0900 265.3000 ;
      RECT 153.8250 19.5000 158.8250 265.3000 ;
      RECT 135.5600 19.5000 150.8250 265.3000 ;
      RECT 127.5600 19.5000 132.5600 265.3000 ;
      RECT 109.2950 19.5000 124.5600 265.3000 ;
      RECT 101.2950 19.5000 106.2950 265.3000 ;
      RECT 83.0300 19.5000 98.2950 265.3000 ;
      RECT 75.0300 19.5000 80.0300 265.3000 ;
      RECT 56.7650 19.5000 72.0300 265.3000 ;
      RECT 48.7650 19.5000 53.7650 265.3000 ;
      RECT 30.5000 19.5000 45.7650 265.3000 ;
      RECT 22.5000 19.5000 27.5000 265.3000 ;
      RECT 258.8850 19.3350 286.4000 19.5000 ;
      RECT 232.6200 19.3350 255.8850 19.5000 ;
      RECT 206.3550 19.3350 229.6200 19.5000 ;
      RECT 180.0900 19.3350 203.3550 19.5000 ;
      RECT 153.8250 19.3350 177.0900 19.5000 ;
      RECT 127.5600 19.3350 150.8250 19.5000 ;
      RECT 101.2950 19.3350 124.5600 19.5000 ;
      RECT 75.0300 19.3350 98.2950 19.5000 ;
      RECT 48.7650 19.3350 72.0300 19.5000 ;
      RECT 22.5000 19.3350 45.7650 19.5000 ;
      RECT 0.0000 19.3350 19.5000 265.4650 ;
      RECT 0.0000 0.0000 286.4000 19.3350 ;
  END
END sram_w16

END LIBRARY
